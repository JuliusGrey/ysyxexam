module iFetch(
  input         clock,
  input         reset,
  input  [31:0] io_instIn,
  output [31:0] io_instOut,
  output [31:0] io_pc,
  output [31:0] io_snpc,
  input  [31:0] io_dnpc,
  input         io_jump,
  input         intrTimeCnt_0,
  input         hazardPCBlock_0,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[Reg.scala 27:20]
  wire [31:0] snpc = pc + 32'h4; // @[iFetch.scala 37:14]
  wire  _T_1 = block1_0 | block23_0; // @[iFetch.scala 35:78]
  wire  _T_2 = ~_T_1; // @[iFetch.scala 35:70]
  wire  _T_3 = ~hazardPCBlock_0; // @[iFetch.scala 35:95]
  wire  _T_4 = _T_3 | intrTimeCnt_0; // @[iFetch.scala 35:110]
  wire  _T_5 = _T_2 & _T_4; // @[iFetch.scala 35:91]
  assign io_instOut = io_instIn; // @[iFetch.scala 52:14]
  assign io_pc = pc; // @[iFetch.scala 45:9]
  assign io_snpc = pc + 32'h4; // @[iFetch.scala 38:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h80000000;
    end else if (_T_5) begin
      if (io_jump) begin
        pc <= io_dnpc;
      end else begin
        pc <= snpc;
      end
    end
  end
endmodule
module immeGen(
  input  [31:0] io_inst,
  output [63:0] io_imme
);
  wire [51:0] _T_3 = io_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Iimm = {_T_3,io_inst[31:20]}; // @[Cat.scala 29:58]
  wire [11:0] _T_6 = {io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 29:58]
  wire [51:0] _T_9 = _T_6[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Simm = {_T_9,io_inst[31:25],io_inst[11:7]}; // @[Cat.scala 29:58]
  wire [12:0] _T_17 = {io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [50:0] _T_20 = _T_17[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Bimm = {_T_20,io_inst[31],io_inst[7],io_inst[30:25],io_inst[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_22 = {io_inst[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_25 = _T_22[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Uimm = {_T_25,io_inst[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [20:0] _T_33 = {io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [42:0] _T_36 = _T_33[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Jimm = {_T_36,io_inst[31],io_inst[19:12],io_inst[20],io_inst[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_37 = io_inst & 32'h707f; // @[immeGen.scala 55:47]
  wire  _T_38 = 32'h1063 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_40 = 32'h23 == _T_37; // @[immeGen.scala 54:47]
  wire  _T_42 = 32'h6003 == _T_37; // @[immeGen.scala 51:47]
  wire [31:0] _T_43 = io_inst & 32'hfc00707f; // @[immeGen.scala 51:47]
  wire  _T_44 = 32'h1013 == _T_43; // @[immeGen.scala 51:47]
  wire  _T_46 = 32'h5003 == _T_37; // @[immeGen.scala 51:47]
  wire [31:0] _T_47 = io_inst & 32'h7f; // @[immeGen.scala 53:47]
  wire  _T_48 = 32'h17 == _T_47; // @[immeGen.scala 53:47]
  wire  _T_50 = 32'h1b == _T_37; // @[immeGen.scala 51:47]
  wire  _T_52 = 32'h3 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_54 = 32'h5063 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_56 = 32'h2023 == _T_37; // @[immeGen.scala 54:47]
  wire  _T_58 = 32'h4003 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_60 = 32'h2003 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_62 = 32'h6f == _T_47; // @[immeGen.scala 52:47]
  wire [31:0] _T_63 = io_inst & 32'hfe00707f; // @[immeGen.scala 51:47]
  wire  _T_64 = 32'h4000501b == _T_63; // @[immeGen.scala 51:47]
  wire  _T_66 = 32'h67 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_68 = 32'h6063 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_70 = 32'h3023 == _T_37; // @[immeGen.scala 54:47]
  wire  _T_72 = 32'h5013 == _T_43; // @[immeGen.scala 51:47]
  wire  _T_74 = 32'h4063 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_76 = 32'h101b == _T_63; // @[immeGen.scala 51:47]
  wire  _T_78 = 32'h37 == _T_47; // @[immeGen.scala 53:47]
  wire  _T_80 = 32'h1023 == _T_37; // @[immeGen.scala 54:47]
  wire  _T_82 = 32'h4013 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_84 = 32'h3013 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_86 = 32'h1003 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_88 = 32'h40005013 == _T_43; // @[immeGen.scala 51:47]
  wire  _T_90 = 32'h3003 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_92 = 32'h13 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_94 = 32'h501b == _T_63; // @[immeGen.scala 51:47]
  wire  _T_96 = 32'h7063 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_98 = 32'h7013 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_100 = 32'h63 == _T_37; // @[immeGen.scala 55:47]
  wire  _T_102 = 32'h6013 == _T_37; // @[immeGen.scala 51:47]
  wire  _T_104 = 32'h1073 == _T_37; // @[immeGen.scala 61:29]
  wire  _T_106 = 32'h2073 == _T_37; // @[immeGen.scala 62:29]
  wire  _T_108 = 32'h6073 == _T_37; // @[immeGen.scala 63:29]
  wire  _T_110 = 32'h7073 == _T_37; // @[immeGen.scala 64:29]
  wire  _T_112 = 32'h3073 == _T_37; // @[immeGen.scala 65:29]
  wire [63:0] _T_113 = _T_112 ? Iimm : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _T_114 = _T_110 ? Iimm : _T_113; // @[Mux.scala 98:16]
  wire [63:0] _T_115 = _T_108 ? Iimm : _T_114; // @[Mux.scala 98:16]
  wire [63:0] _T_116 = _T_106 ? Iimm : _T_115; // @[Mux.scala 98:16]
  wire [63:0] _T_117 = _T_104 ? Iimm : _T_116; // @[Mux.scala 98:16]
  wire [63:0] _T_118 = _T_102 ? Iimm : _T_117; // @[Mux.scala 98:16]
  wire [63:0] _T_119 = _T_100 ? Bimm : _T_118; // @[Mux.scala 98:16]
  wire [63:0] _T_120 = _T_98 ? Iimm : _T_119; // @[Mux.scala 98:16]
  wire [63:0] _T_121 = _T_96 ? Bimm : _T_120; // @[Mux.scala 98:16]
  wire [63:0] _T_122 = _T_94 ? Iimm : _T_121; // @[Mux.scala 98:16]
  wire [63:0] _T_123 = _T_92 ? Iimm : _T_122; // @[Mux.scala 98:16]
  wire [63:0] _T_124 = _T_90 ? Iimm : _T_123; // @[Mux.scala 98:16]
  wire [63:0] _T_125 = _T_88 ? Iimm : _T_124; // @[Mux.scala 98:16]
  wire [63:0] _T_126 = _T_86 ? Iimm : _T_125; // @[Mux.scala 98:16]
  wire [63:0] _T_127 = _T_84 ? Iimm : _T_126; // @[Mux.scala 98:16]
  wire [63:0] _T_128 = _T_82 ? Iimm : _T_127; // @[Mux.scala 98:16]
  wire [63:0] _T_129 = _T_80 ? Simm : _T_128; // @[Mux.scala 98:16]
  wire [63:0] _T_130 = _T_78 ? Uimm : _T_129; // @[Mux.scala 98:16]
  wire [63:0] _T_131 = _T_76 ? Iimm : _T_130; // @[Mux.scala 98:16]
  wire [63:0] _T_132 = _T_74 ? Bimm : _T_131; // @[Mux.scala 98:16]
  wire [63:0] _T_133 = _T_72 ? Iimm : _T_132; // @[Mux.scala 98:16]
  wire [63:0] _T_134 = _T_70 ? Simm : _T_133; // @[Mux.scala 98:16]
  wire [63:0] _T_135 = _T_68 ? Bimm : _T_134; // @[Mux.scala 98:16]
  wire [63:0] _T_136 = _T_66 ? Iimm : _T_135; // @[Mux.scala 98:16]
  wire [63:0] _T_137 = _T_64 ? Iimm : _T_136; // @[Mux.scala 98:16]
  wire [63:0] _T_138 = _T_62 ? Jimm : _T_137; // @[Mux.scala 98:16]
  wire [63:0] _T_139 = _T_60 ? Iimm : _T_138; // @[Mux.scala 98:16]
  wire [63:0] _T_140 = _T_58 ? Iimm : _T_139; // @[Mux.scala 98:16]
  wire [63:0] _T_141 = _T_56 ? Simm : _T_140; // @[Mux.scala 98:16]
  wire [63:0] _T_142 = _T_54 ? Bimm : _T_141; // @[Mux.scala 98:16]
  wire [63:0] _T_143 = _T_52 ? Iimm : _T_142; // @[Mux.scala 98:16]
  wire [63:0] _T_144 = _T_50 ? Iimm : _T_143; // @[Mux.scala 98:16]
  wire [63:0] _T_145 = _T_48 ? Uimm : _T_144; // @[Mux.scala 98:16]
  wire [63:0] _T_146 = _T_46 ? Iimm : _T_145; // @[Mux.scala 98:16]
  wire [63:0] _T_147 = _T_44 ? Iimm : _T_146; // @[Mux.scala 98:16]
  wire [63:0] _T_148 = _T_42 ? Iimm : _T_147; // @[Mux.scala 98:16]
  wire [63:0] _T_149 = _T_40 ? Simm : _T_148; // @[Mux.scala 98:16]
  assign io_imme = _T_38 ? Bimm : _T_149; // @[immeGen.scala 67:13]
endmodule
module RF(
  input         clock,
  input  [31:0] io_pc,
  input         io_we,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  output [63:0] io_dout1,
  output [63:0] io_dout2,
  input  [63:0] io_din,
  input  [4:0]  io_rsWB,
  output [63:0] io_doutWB,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] DPIC_RegRead_ins_inst_0; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_1; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_2; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_3; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_4; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_5; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_6; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_7; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_8; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_9; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_10; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_11; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_12; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_13; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_14; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_15; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_16; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_17; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_18; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_19; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_20; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_21; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_22; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_23; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_24; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_25; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_26; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_27; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_28; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_29; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_30; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_inst_31; // @[regFile.scala 27:32]
  wire [63:0] DPIC_RegRead_ins_pc; // @[regFile.scala 27:32]
  wire  _T_1 = block1_0 | block23_0; // @[regFile.scala 61:50]
  wire  _T_2 = ~_T_1; // @[regFile.scala 61:41]
  wire  _T_6 = io_rd == 5'h1; // @[regFile.scala 49:22]
  wire  _T_7 = io_we & _T_6; // @[regFile.scala 49:13]
  wire  _T_10 = _T_7 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_11; // @[Reg.scala 15:16]
  wire  _T_13 = io_rd == 5'h2; // @[regFile.scala 49:22]
  wire  _T_14 = io_we & _T_13; // @[regFile.scala 49:13]
  wire  _T_17 = _T_14 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_18; // @[Reg.scala 15:16]
  wire  _T_20 = io_rd == 5'h3; // @[regFile.scala 49:22]
  wire  _T_21 = io_we & _T_20; // @[regFile.scala 49:13]
  wire  _T_24 = _T_21 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_25; // @[Reg.scala 15:16]
  wire  _T_27 = io_rd == 5'h4; // @[regFile.scala 49:22]
  wire  _T_28 = io_we & _T_27; // @[regFile.scala 49:13]
  wire  _T_31 = _T_28 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_32; // @[Reg.scala 15:16]
  wire  _T_34 = io_rd == 5'h5; // @[regFile.scala 49:22]
  wire  _T_35 = io_we & _T_34; // @[regFile.scala 49:13]
  wire  _T_38 = _T_35 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_39; // @[Reg.scala 15:16]
  wire  _T_41 = io_rd == 5'h6; // @[regFile.scala 49:22]
  wire  _T_42 = io_we & _T_41; // @[regFile.scala 49:13]
  wire  _T_45 = _T_42 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_46; // @[Reg.scala 15:16]
  wire  _T_48 = io_rd == 5'h7; // @[regFile.scala 49:22]
  wire  _T_49 = io_we & _T_48; // @[regFile.scala 49:13]
  wire  _T_52 = _T_49 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_53; // @[Reg.scala 15:16]
  wire  _T_55 = io_rd == 5'h8; // @[regFile.scala 49:22]
  wire  _T_56 = io_we & _T_55; // @[regFile.scala 49:13]
  wire  _T_59 = _T_56 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_60; // @[Reg.scala 15:16]
  wire  _T_62 = io_rd == 5'h9; // @[regFile.scala 49:22]
  wire  _T_63 = io_we & _T_62; // @[regFile.scala 49:13]
  wire  _T_66 = _T_63 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_67; // @[Reg.scala 15:16]
  wire  _T_69 = io_rd == 5'ha; // @[regFile.scala 49:22]
  wire  _T_70 = io_we & _T_69; // @[regFile.scala 49:13]
  wire  _T_73 = _T_70 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_74; // @[Reg.scala 15:16]
  wire  _T_76 = io_rd == 5'hb; // @[regFile.scala 49:22]
  wire  _T_77 = io_we & _T_76; // @[regFile.scala 49:13]
  wire  _T_80 = _T_77 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_81; // @[Reg.scala 15:16]
  wire  _T_83 = io_rd == 5'hc; // @[regFile.scala 49:22]
  wire  _T_84 = io_we & _T_83; // @[regFile.scala 49:13]
  wire  _T_87 = _T_84 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_88; // @[Reg.scala 15:16]
  wire  _T_90 = io_rd == 5'hd; // @[regFile.scala 49:22]
  wire  _T_91 = io_we & _T_90; // @[regFile.scala 49:13]
  wire  _T_94 = _T_91 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_95; // @[Reg.scala 15:16]
  wire  _T_97 = io_rd == 5'he; // @[regFile.scala 49:22]
  wire  _T_98 = io_we & _T_97; // @[regFile.scala 49:13]
  wire  _T_101 = _T_98 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_102; // @[Reg.scala 15:16]
  wire  _T_104 = io_rd == 5'hf; // @[regFile.scala 49:22]
  wire  _T_105 = io_we & _T_104; // @[regFile.scala 49:13]
  wire  _T_108 = _T_105 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_109; // @[Reg.scala 15:16]
  wire  _T_111 = io_rd == 5'h10; // @[regFile.scala 49:22]
  wire  _T_112 = io_we & _T_111; // @[regFile.scala 49:13]
  wire  _T_115 = _T_112 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_116; // @[Reg.scala 15:16]
  wire  _T_118 = io_rd == 5'h11; // @[regFile.scala 49:22]
  wire  _T_119 = io_we & _T_118; // @[regFile.scala 49:13]
  wire  _T_122 = _T_119 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_123; // @[Reg.scala 15:16]
  wire  _T_125 = io_rd == 5'h12; // @[regFile.scala 49:22]
  wire  _T_126 = io_we & _T_125; // @[regFile.scala 49:13]
  wire  _T_129 = _T_126 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_130; // @[Reg.scala 15:16]
  wire  _T_132 = io_rd == 5'h13; // @[regFile.scala 49:22]
  wire  _T_133 = io_we & _T_132; // @[regFile.scala 49:13]
  wire  _T_136 = _T_133 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_137; // @[Reg.scala 15:16]
  wire  _T_139 = io_rd == 5'h14; // @[regFile.scala 49:22]
  wire  _T_140 = io_we & _T_139; // @[regFile.scala 49:13]
  wire  _T_143 = _T_140 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_144; // @[Reg.scala 15:16]
  wire  _T_146 = io_rd == 5'h15; // @[regFile.scala 49:22]
  wire  _T_147 = io_we & _T_146; // @[regFile.scala 49:13]
  wire  _T_150 = _T_147 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_151; // @[Reg.scala 15:16]
  wire  _T_153 = io_rd == 5'h16; // @[regFile.scala 49:22]
  wire  _T_154 = io_we & _T_153; // @[regFile.scala 49:13]
  wire  _T_157 = _T_154 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_158; // @[Reg.scala 15:16]
  wire  _T_160 = io_rd == 5'h17; // @[regFile.scala 49:22]
  wire  _T_161 = io_we & _T_160; // @[regFile.scala 49:13]
  wire  _T_164 = _T_161 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_165; // @[Reg.scala 15:16]
  wire  _T_167 = io_rd == 5'h18; // @[regFile.scala 49:22]
  wire  _T_168 = io_we & _T_167; // @[regFile.scala 49:13]
  wire  _T_171 = _T_168 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_172; // @[Reg.scala 15:16]
  wire  _T_174 = io_rd == 5'h19; // @[regFile.scala 49:22]
  wire  _T_175 = io_we & _T_174; // @[regFile.scala 49:13]
  wire  _T_178 = _T_175 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_179; // @[Reg.scala 15:16]
  wire  _T_181 = io_rd == 5'h1a; // @[regFile.scala 49:22]
  wire  _T_182 = io_we & _T_181; // @[regFile.scala 49:13]
  wire  _T_185 = _T_182 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_186; // @[Reg.scala 15:16]
  wire  _T_188 = io_rd == 5'h1b; // @[regFile.scala 49:22]
  wire  _T_189 = io_we & _T_188; // @[regFile.scala 49:13]
  wire  _T_192 = _T_189 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_193; // @[Reg.scala 15:16]
  wire  _T_195 = io_rd == 5'h1c; // @[regFile.scala 49:22]
  wire  _T_196 = io_we & _T_195; // @[regFile.scala 49:13]
  wire  _T_199 = _T_196 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_200; // @[Reg.scala 15:16]
  wire  _T_202 = io_rd == 5'h1d; // @[regFile.scala 49:22]
  wire  _T_203 = io_we & _T_202; // @[regFile.scala 49:13]
  wire  _T_206 = _T_203 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_207; // @[Reg.scala 15:16]
  wire  _T_209 = io_rd == 5'h1e; // @[regFile.scala 49:22]
  wire  _T_210 = io_we & _T_209; // @[regFile.scala 49:13]
  wire  _T_213 = _T_210 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_214; // @[Reg.scala 15:16]
  wire  _T_216 = io_rd == 5'h1f; // @[regFile.scala 49:22]
  wire  _T_217 = io_we & _T_216; // @[regFile.scala 49:13]
  wire  _T_220 = _T_217 & _T_2; // @[regFile.scala 61:38]
  reg [63:0] _T_221; // @[Reg.scala 15:16]
  wire  _T_222 = 5'h1 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_223 = _T_222 ? _T_11 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_224 = 5'h2 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_225 = _T_224 ? _T_18 : _T_223; // @[Mux.scala 80:57]
  wire  _T_226 = 5'h3 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_227 = _T_226 ? _T_25 : _T_225; // @[Mux.scala 80:57]
  wire  _T_228 = 5'h4 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_229 = _T_228 ? _T_32 : _T_227; // @[Mux.scala 80:57]
  wire  _T_230 = 5'h5 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_231 = _T_230 ? _T_39 : _T_229; // @[Mux.scala 80:57]
  wire  _T_232 = 5'h6 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_233 = _T_232 ? _T_46 : _T_231; // @[Mux.scala 80:57]
  wire  _T_234 = 5'h7 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_235 = _T_234 ? _T_53 : _T_233; // @[Mux.scala 80:57]
  wire  _T_236 = 5'h8 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_237 = _T_236 ? _T_60 : _T_235; // @[Mux.scala 80:57]
  wire  _T_238 = 5'h9 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_239 = _T_238 ? _T_67 : _T_237; // @[Mux.scala 80:57]
  wire  _T_240 = 5'ha == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_241 = _T_240 ? _T_74 : _T_239; // @[Mux.scala 80:57]
  wire  _T_242 = 5'hb == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_243 = _T_242 ? _T_81 : _T_241; // @[Mux.scala 80:57]
  wire  _T_244 = 5'hc == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_245 = _T_244 ? _T_88 : _T_243; // @[Mux.scala 80:57]
  wire  _T_246 = 5'hd == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_247 = _T_246 ? _T_95 : _T_245; // @[Mux.scala 80:57]
  wire  _T_248 = 5'he == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_249 = _T_248 ? _T_102 : _T_247; // @[Mux.scala 80:57]
  wire  _T_250 = 5'hf == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_251 = _T_250 ? _T_109 : _T_249; // @[Mux.scala 80:57]
  wire  _T_252 = 5'h10 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_253 = _T_252 ? _T_116 : _T_251; // @[Mux.scala 80:57]
  wire  _T_254 = 5'h11 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_255 = _T_254 ? _T_123 : _T_253; // @[Mux.scala 80:57]
  wire  _T_256 = 5'h12 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_257 = _T_256 ? _T_130 : _T_255; // @[Mux.scala 80:57]
  wire  _T_258 = 5'h13 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_259 = _T_258 ? _T_137 : _T_257; // @[Mux.scala 80:57]
  wire  _T_260 = 5'h14 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_261 = _T_260 ? _T_144 : _T_259; // @[Mux.scala 80:57]
  wire  _T_262 = 5'h15 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_263 = _T_262 ? _T_151 : _T_261; // @[Mux.scala 80:57]
  wire  _T_264 = 5'h16 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_265 = _T_264 ? _T_158 : _T_263; // @[Mux.scala 80:57]
  wire  _T_266 = 5'h17 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_267 = _T_266 ? _T_165 : _T_265; // @[Mux.scala 80:57]
  wire  _T_268 = 5'h18 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_269 = _T_268 ? _T_172 : _T_267; // @[Mux.scala 80:57]
  wire  _T_270 = 5'h19 == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_271 = _T_270 ? _T_179 : _T_269; // @[Mux.scala 80:57]
  wire  _T_272 = 5'h1a == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_273 = _T_272 ? _T_186 : _T_271; // @[Mux.scala 80:57]
  wire  _T_274 = 5'h1b == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_275 = _T_274 ? _T_193 : _T_273; // @[Mux.scala 80:57]
  wire  _T_276 = 5'h1c == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_277 = _T_276 ? _T_200 : _T_275; // @[Mux.scala 80:57]
  wire  _T_278 = 5'h1d == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_279 = _T_278 ? _T_207 : _T_277; // @[Mux.scala 80:57]
  wire  _T_280 = 5'h1e == io_rs1; // @[Mux.scala 80:60]
  wire [63:0] _T_281 = _T_280 ? _T_214 : _T_279; // @[Mux.scala 80:57]
  wire  _T_282 = 5'h1f == io_rs1; // @[Mux.scala 80:60]
  wire  _T_284 = 5'h1 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_285 = _T_284 ? _T_11 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_286 = 5'h2 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_287 = _T_286 ? _T_18 : _T_285; // @[Mux.scala 80:57]
  wire  _T_288 = 5'h3 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_289 = _T_288 ? _T_25 : _T_287; // @[Mux.scala 80:57]
  wire  _T_290 = 5'h4 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_291 = _T_290 ? _T_32 : _T_289; // @[Mux.scala 80:57]
  wire  _T_292 = 5'h5 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_293 = _T_292 ? _T_39 : _T_291; // @[Mux.scala 80:57]
  wire  _T_294 = 5'h6 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_295 = _T_294 ? _T_46 : _T_293; // @[Mux.scala 80:57]
  wire  _T_296 = 5'h7 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_297 = _T_296 ? _T_53 : _T_295; // @[Mux.scala 80:57]
  wire  _T_298 = 5'h8 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_299 = _T_298 ? _T_60 : _T_297; // @[Mux.scala 80:57]
  wire  _T_300 = 5'h9 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_301 = _T_300 ? _T_67 : _T_299; // @[Mux.scala 80:57]
  wire  _T_302 = 5'ha == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_303 = _T_302 ? _T_74 : _T_301; // @[Mux.scala 80:57]
  wire  _T_304 = 5'hb == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_305 = _T_304 ? _T_81 : _T_303; // @[Mux.scala 80:57]
  wire  _T_306 = 5'hc == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_307 = _T_306 ? _T_88 : _T_305; // @[Mux.scala 80:57]
  wire  _T_308 = 5'hd == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_309 = _T_308 ? _T_95 : _T_307; // @[Mux.scala 80:57]
  wire  _T_310 = 5'he == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_311 = _T_310 ? _T_102 : _T_309; // @[Mux.scala 80:57]
  wire  _T_312 = 5'hf == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_313 = _T_312 ? _T_109 : _T_311; // @[Mux.scala 80:57]
  wire  _T_314 = 5'h10 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_315 = _T_314 ? _T_116 : _T_313; // @[Mux.scala 80:57]
  wire  _T_316 = 5'h11 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_317 = _T_316 ? _T_123 : _T_315; // @[Mux.scala 80:57]
  wire  _T_318 = 5'h12 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_319 = _T_318 ? _T_130 : _T_317; // @[Mux.scala 80:57]
  wire  _T_320 = 5'h13 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_321 = _T_320 ? _T_137 : _T_319; // @[Mux.scala 80:57]
  wire  _T_322 = 5'h14 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_323 = _T_322 ? _T_144 : _T_321; // @[Mux.scala 80:57]
  wire  _T_324 = 5'h15 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_325 = _T_324 ? _T_151 : _T_323; // @[Mux.scala 80:57]
  wire  _T_326 = 5'h16 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_327 = _T_326 ? _T_158 : _T_325; // @[Mux.scala 80:57]
  wire  _T_328 = 5'h17 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_329 = _T_328 ? _T_165 : _T_327; // @[Mux.scala 80:57]
  wire  _T_330 = 5'h18 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_331 = _T_330 ? _T_172 : _T_329; // @[Mux.scala 80:57]
  wire  _T_332 = 5'h19 == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_333 = _T_332 ? _T_179 : _T_331; // @[Mux.scala 80:57]
  wire  _T_334 = 5'h1a == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_335 = _T_334 ? _T_186 : _T_333; // @[Mux.scala 80:57]
  wire  _T_336 = 5'h1b == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_337 = _T_336 ? _T_193 : _T_335; // @[Mux.scala 80:57]
  wire  _T_338 = 5'h1c == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_339 = _T_338 ? _T_200 : _T_337; // @[Mux.scala 80:57]
  wire  _T_340 = 5'h1d == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_341 = _T_340 ? _T_207 : _T_339; // @[Mux.scala 80:57]
  wire  _T_342 = 5'h1e == io_rs2; // @[Mux.scala 80:60]
  wire [63:0] _T_343 = _T_342 ? _T_214 : _T_341; // @[Mux.scala 80:57]
  wire  _T_344 = 5'h1f == io_rs2; // @[Mux.scala 80:60]
  wire  _T_346 = 5'h1 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_347 = _T_346 ? _T_11 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_348 = 5'h2 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_349 = _T_348 ? _T_18 : _T_347; // @[Mux.scala 80:57]
  wire  _T_350 = 5'h3 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_351 = _T_350 ? _T_25 : _T_349; // @[Mux.scala 80:57]
  wire  _T_352 = 5'h4 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_353 = _T_352 ? _T_32 : _T_351; // @[Mux.scala 80:57]
  wire  _T_354 = 5'h5 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_355 = _T_354 ? _T_39 : _T_353; // @[Mux.scala 80:57]
  wire  _T_356 = 5'h6 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_357 = _T_356 ? _T_46 : _T_355; // @[Mux.scala 80:57]
  wire  _T_358 = 5'h7 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_359 = _T_358 ? _T_53 : _T_357; // @[Mux.scala 80:57]
  wire  _T_360 = 5'h8 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_361 = _T_360 ? _T_60 : _T_359; // @[Mux.scala 80:57]
  wire  _T_362 = 5'h9 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_363 = _T_362 ? _T_67 : _T_361; // @[Mux.scala 80:57]
  wire  _T_364 = 5'ha == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_365 = _T_364 ? _T_74 : _T_363; // @[Mux.scala 80:57]
  wire  _T_366 = 5'hb == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_367 = _T_366 ? _T_81 : _T_365; // @[Mux.scala 80:57]
  wire  _T_368 = 5'hc == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_369 = _T_368 ? _T_88 : _T_367; // @[Mux.scala 80:57]
  wire  _T_370 = 5'hd == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_371 = _T_370 ? _T_95 : _T_369; // @[Mux.scala 80:57]
  wire  _T_372 = 5'he == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_373 = _T_372 ? _T_102 : _T_371; // @[Mux.scala 80:57]
  wire  _T_374 = 5'hf == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_375 = _T_374 ? _T_109 : _T_373; // @[Mux.scala 80:57]
  wire  _T_376 = 5'h10 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_377 = _T_376 ? _T_116 : _T_375; // @[Mux.scala 80:57]
  wire  _T_378 = 5'h11 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_379 = _T_378 ? _T_123 : _T_377; // @[Mux.scala 80:57]
  wire  _T_380 = 5'h12 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_381 = _T_380 ? _T_130 : _T_379; // @[Mux.scala 80:57]
  wire  _T_382 = 5'h13 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_383 = _T_382 ? _T_137 : _T_381; // @[Mux.scala 80:57]
  wire  _T_384 = 5'h14 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_385 = _T_384 ? _T_144 : _T_383; // @[Mux.scala 80:57]
  wire  _T_386 = 5'h15 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_387 = _T_386 ? _T_151 : _T_385; // @[Mux.scala 80:57]
  wire  _T_388 = 5'h16 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_389 = _T_388 ? _T_158 : _T_387; // @[Mux.scala 80:57]
  wire  _T_390 = 5'h17 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_391 = _T_390 ? _T_165 : _T_389; // @[Mux.scala 80:57]
  wire  _T_392 = 5'h18 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_393 = _T_392 ? _T_172 : _T_391; // @[Mux.scala 80:57]
  wire  _T_394 = 5'h19 == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_395 = _T_394 ? _T_179 : _T_393; // @[Mux.scala 80:57]
  wire  _T_396 = 5'h1a == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_397 = _T_396 ? _T_186 : _T_395; // @[Mux.scala 80:57]
  wire  _T_398 = 5'h1b == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_399 = _T_398 ? _T_193 : _T_397; // @[Mux.scala 80:57]
  wire  _T_400 = 5'h1c == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_401 = _T_400 ? _T_200 : _T_399; // @[Mux.scala 80:57]
  wire  _T_402 = 5'h1d == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_403 = _T_402 ? _T_207 : _T_401; // @[Mux.scala 80:57]
  wire  _T_404 = 5'h1e == io_rsWB; // @[Mux.scala 80:60]
  wire [63:0] _T_405 = _T_404 ? _T_214 : _T_403; // @[Mux.scala 80:57]
  wire  _T_406 = 5'h1f == io_rsWB; // @[Mux.scala 80:60]
  DPIC_RegRead DPIC_RegRead_ins ( // @[regFile.scala 27:32]
    .inst_0(DPIC_RegRead_ins_inst_0),
    .inst_1(DPIC_RegRead_ins_inst_1),
    .inst_2(DPIC_RegRead_ins_inst_2),
    .inst_3(DPIC_RegRead_ins_inst_3),
    .inst_4(DPIC_RegRead_ins_inst_4),
    .inst_5(DPIC_RegRead_ins_inst_5),
    .inst_6(DPIC_RegRead_ins_inst_6),
    .inst_7(DPIC_RegRead_ins_inst_7),
    .inst_8(DPIC_RegRead_ins_inst_8),
    .inst_9(DPIC_RegRead_ins_inst_9),
    .inst_10(DPIC_RegRead_ins_inst_10),
    .inst_11(DPIC_RegRead_ins_inst_11),
    .inst_12(DPIC_RegRead_ins_inst_12),
    .inst_13(DPIC_RegRead_ins_inst_13),
    .inst_14(DPIC_RegRead_ins_inst_14),
    .inst_15(DPIC_RegRead_ins_inst_15),
    .inst_16(DPIC_RegRead_ins_inst_16),
    .inst_17(DPIC_RegRead_ins_inst_17),
    .inst_18(DPIC_RegRead_ins_inst_18),
    .inst_19(DPIC_RegRead_ins_inst_19),
    .inst_20(DPIC_RegRead_ins_inst_20),
    .inst_21(DPIC_RegRead_ins_inst_21),
    .inst_22(DPIC_RegRead_ins_inst_22),
    .inst_23(DPIC_RegRead_ins_inst_23),
    .inst_24(DPIC_RegRead_ins_inst_24),
    .inst_25(DPIC_RegRead_ins_inst_25),
    .inst_26(DPIC_RegRead_ins_inst_26),
    .inst_27(DPIC_RegRead_ins_inst_27),
    .inst_28(DPIC_RegRead_ins_inst_28),
    .inst_29(DPIC_RegRead_ins_inst_29),
    .inst_30(DPIC_RegRead_ins_inst_30),
    .inst_31(DPIC_RegRead_ins_inst_31),
    .pc(DPIC_RegRead_ins_pc)
  );
  assign io_dout1 = _T_282 ? _T_221 : _T_281; // @[regFile.scala 66:12]
  assign io_dout2 = _T_344 ? _T_221 : _T_343; // @[regFile.scala 67:12]
  assign io_doutWB = _T_406 ? _T_221 : _T_405; // @[regFile.scala 69:13]
  assign DPIC_RegRead_ins_inst_0 = 64'h0; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_1 = _T_11; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_2 = _T_18; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_3 = _T_25; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_4 = _T_32; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_5 = _T_39; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_6 = _T_46; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_7 = _T_53; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_8 = _T_60; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_9 = _T_67; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_10 = _T_74; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_11 = _T_81; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_12 = _T_88; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_13 = _T_95; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_14 = _T_102; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_15 = _T_109; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_16 = _T_116; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_17 = _T_123; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_18 = _T_130; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_19 = _T_137; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_20 = _T_144; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_21 = _T_151; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_22 = _T_158; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_23 = _T_165; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_24 = _T_172; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_25 = _T_179; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_26 = _T_186; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_27 = _T_193; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_28 = _T_200; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_29 = _T_207; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_30 = _T_214; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_inst_31 = _T_221; // @[regFile.scala 62:33]
  assign DPIC_RegRead_ins_pc = {{32'd0}, io_pc}; // @[regFile.scala 28:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_11 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_18 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_25 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_32 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  _T_46 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  _T_53 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_60 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_67 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_74 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  _T_81 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  _T_88 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  _T_95 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  _T_102 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  _T_109 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  _T_116 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  _T_123 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  _T_130 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  _T_137 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_144 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_151 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_158 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  _T_165 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_172 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_179 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_186 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_193 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_200 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  _T_207 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  _T_214 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_221 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T_11 <= io_din;
    end
    if (_T_17) begin
      _T_18 <= io_din;
    end
    if (_T_24) begin
      _T_25 <= io_din;
    end
    if (_T_31) begin
      _T_32 <= io_din;
    end
    if (_T_38) begin
      _T_39 <= io_din;
    end
    if (_T_45) begin
      _T_46 <= io_din;
    end
    if (_T_52) begin
      _T_53 <= io_din;
    end
    if (_T_59) begin
      _T_60 <= io_din;
    end
    if (_T_66) begin
      _T_67 <= io_din;
    end
    if (_T_73) begin
      _T_74 <= io_din;
    end
    if (_T_80) begin
      _T_81 <= io_din;
    end
    if (_T_87) begin
      _T_88 <= io_din;
    end
    if (_T_94) begin
      _T_95 <= io_din;
    end
    if (_T_101) begin
      _T_102 <= io_din;
    end
    if (_T_108) begin
      _T_109 <= io_din;
    end
    if (_T_115) begin
      _T_116 <= io_din;
    end
    if (_T_122) begin
      _T_123 <= io_din;
    end
    if (_T_129) begin
      _T_130 <= io_din;
    end
    if (_T_136) begin
      _T_137 <= io_din;
    end
    if (_T_143) begin
      _T_144 <= io_din;
    end
    if (_T_150) begin
      _T_151 <= io_din;
    end
    if (_T_157) begin
      _T_158 <= io_din;
    end
    if (_T_164) begin
      _T_165 <= io_din;
    end
    if (_T_171) begin
      _T_172 <= io_din;
    end
    if (_T_178) begin
      _T_179 <= io_din;
    end
    if (_T_185) begin
      _T_186 <= io_din;
    end
    if (_T_192) begin
      _T_193 <= io_din;
    end
    if (_T_199) begin
      _T_200 <= io_din;
    end
    if (_T_206) begin
      _T_207 <= io_din;
    end
    if (_T_213) begin
      _T_214 <= io_din;
    end
    if (_T_220) begin
      _T_221 <= io_din;
    end
  end
endmodule
module iDecode(
  input         clock,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_regEn,
  output [63:0] io_dataEx_imme,
  output [63:0] io_dataEx_dOut1,
  output [63:0] io_dataEx_dOut2,
  input  [63:0] io_dataEx_dIn,
  output [4:0]  io_rdOut,
  input  [4:0]  io_rdIn,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  input  [4:0]  io_rsWB,
  output [63:0] io_dOutWB,
  input         block1,
  input         block23
);
  wire [31:0] imme_io_inst; // @[iDecode.scala 28:19]
  wire [63:0] imme_io_imme; // @[iDecode.scala 28:19]
  wire  rf_clock; // @[iDecode.scala 42:18]
  wire [31:0] rf_io_pc; // @[iDecode.scala 42:18]
  wire  rf_io_we; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs1; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs2; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rd; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout1; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout2; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_din; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rsWB; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_doutWB; // @[iDecode.scala 42:18]
  wire  rf_block1_0; // @[iDecode.scala 42:18]
  wire  rf_block23_0; // @[iDecode.scala 42:18]
  immeGen imme ( // @[iDecode.scala 28:19]
    .io_inst(imme_io_inst),
    .io_imme(imme_io_imme)
  );
  RF rf ( // @[iDecode.scala 42:18]
    .clock(rf_clock),
    .io_pc(rf_io_pc),
    .io_we(rf_io_we),
    .io_rs1(rf_io_rs1),
    .io_rs2(rf_io_rs2),
    .io_rd(rf_io_rd),
    .io_dout1(rf_io_dout1),
    .io_dout2(rf_io_dout2),
    .io_din(rf_io_din),
    .io_rsWB(rf_io_rsWB),
    .io_doutWB(rf_io_doutWB),
    .block1_0(rf_block1_0),
    .block23_0(rf_block23_0)
  );
  assign io_dataEx_imme = imme_io_imme; // @[iDecode.scala 30:18]
  assign io_dataEx_dOut1 = rf_io_dout1; // @[iDecode.scala 48:19]
  assign io_dataEx_dOut2 = rf_io_dout2; // @[iDecode.scala 49:19]
  assign io_rdOut = io_inst[11:7]; // @[iDecode.scala 37:12]
  assign io_rs1 = io_inst[19:15]; // @[iDecode.scala 38:10]
  assign io_rs2 = io_inst[24:20]; // @[iDecode.scala 39:10]
  assign io_dOutWB = rf_io_doutWB; // @[iDecode.scala 54:13]
  assign imme_io_inst = io_inst; // @[iDecode.scala 29:16]
  assign rf_clock = clock;
  assign rf_io_pc = io_pc; // @[iDecode.scala 51:12]
  assign rf_io_we = io_regEn; // @[iDecode.scala 46:12]
  assign rf_io_rs1 = io_inst[19:15]; // @[iDecode.scala 43:13]
  assign rf_io_rs2 = io_inst[24:20]; // @[iDecode.scala 44:13]
  assign rf_io_rd = io_rdIn; // @[iDecode.scala 45:12]
  assign rf_io_din = io_dataEx_dIn; // @[iDecode.scala 47:13]
  assign rf_io_rsWB = io_rsWB; // @[iDecode.scala 53:14]
  assign rf_block1_0 = block1;
  assign rf_block23_0 = block23;
endmodule
module add(
  input         io_cin,
  input  [63:0] io_a,
  input  [63:0] io_b,
  output [63:0] io_sum,
  output        io_cout
);
  wire [64:0] _T_1 = {1'h0,io_a}; // @[Cat.scala 29:58]
  wire [64:0] _T_2 = {1'h0,io_b}; // @[Cat.scala 29:58]
  wire [64:0] _T_4 = _T_1 + _T_2; // @[add.scala 17:31]
  wire [64:0] _GEN_0 = {{64'd0}, io_cin}; // @[add.scala 17:52]
  wire [64:0] _T_6 = _T_4 + _GEN_0; // @[add.scala 17:52]
  assign io_sum = _T_6[63:0]; // @[add.scala 18:12]
  assign io_cout = _T_6[64]; // @[add.scala 19:13]
endmodule
module divR2(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_divw,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = io_dividend[63] & io_div_signed; // @[divR2.scala 21:51]
  wire [63:0] _T_2 = ~io_dividend; // @[divR2.scala 21:70]
  wire [63:0] _T_4 = _T_2 + 64'h1; // @[divR2.scala 21:91]
  wire [63:0] dividend64Real = _T_1 ? _T_4 : io_dividend; // @[divR2.scala 21:27]
  wire  _T_6 = io_divisor[63] & io_div_signed; // @[divR2.scala 22:49]
  wire [63:0] _T_7 = ~io_divisor; // @[divR2.scala 22:68]
  wire [63:0] _T_9 = _T_7 + 64'h1; // @[divR2.scala 22:88]
  wire [63:0] divisor64Real = _T_6 ? _T_9 : io_divisor; // @[divR2.scala 22:26]
  wire  _T_12 = io_dividend[63] ^ io_divisor[63]; // @[divR2.scala 23:42]
  wire  quoSgn64 = _T_12 & io_div_signed; // @[divR2.scala 23:67]
  wire  _T_15 = io_dividend[31] & io_div_signed; // @[divR2.scala 26:48]
  wire [31:0] _T_17 = ~io_dividend[31:0]; // @[divR2.scala 26:67]
  wire [31:0] _T_19 = _T_17 + 32'h1; // @[divR2.scala 26:94]
  wire [31:0] dividend32Real = _T_15 ? _T_19 : io_dividend[31:0]; // @[divR2.scala 26:27]
  wire  _T_22 = io_divisor[31] & io_div_signed; // @[divR2.scala 27:46]
  wire [31:0] _T_24 = ~io_divisor[31:0]; // @[divR2.scala 27:65]
  wire [31:0] _T_26 = _T_24 + 32'h1; // @[divR2.scala 27:91]
  wire [31:0] divisor32Real = _T_22 ? _T_26 : io_divisor[31:0]; // @[divR2.scala 27:26]
  wire  _T_30 = io_dividend[31] ^ io_divisor[31]; // @[divR2.scala 28:39]
  wire  quoSgn32 = _T_30 & io_div_signed; // @[divR2.scala 28:61]
  reg [1:0] stateReg; // @[divR2.scala 35:25]
  wire  isDiv32 = stateReg == 2'h1; // @[divR2.scala 37:25]
  wire  isDiv64 = stateReg == 2'h2; // @[divR2.scala 38:26]
  reg [5:0] cnt; // @[divR2.scala 40:20]
  wire [1:0] _T_32 = {io_div_valid,io_divw}; // @[Cat.scala 29:58]
  wire  _T_33 = 2'h3 == _T_32; // @[Mux.scala 80:60]
  wire  _T_35 = 2'h2 == _T_32; // @[Mux.scala 80:60]
  wire  _T_36 = cnt == 6'h1f; // @[divR2.scala 49:26]
  wire  _T_37 = cnt == 6'h3f; // @[divR2.scala 50:26]
  wire  _T_38 = 2'h1 == stateReg; // @[Mux.scala 80:60]
  wire  _T_40 = 2'h2 == stateReg; // @[Mux.scala 80:60]
  wire  _T_42 = 2'h3 == stateReg; // @[Mux.scala 80:60]
  wire  _T_44 = isDiv32 | isDiv64; // @[divR2.scala 63:21]
  wire [5:0] _T_46 = cnt + 6'h1; // @[divR2.scala 63:38]
  reg [127:0] dividendReg; // @[divR2.scala 66:28]
  reg [63:0] resReg; // @[divR2.scala 67:23]
  wire [127:0] _T_51 = {96'h0,dividend32Real}; // @[Cat.scala 29:58]
  wire [127:0] _T_52 = {64'h0,dividend64Real}; // @[Cat.scala 29:58]
  wire [32:0] subed32 = dividendReg[63:31]; // @[divR2.scala 95:27]
  wire [32:0] _GEN_0 = {{1'd0}, divisor32Real}; // @[divR2.scala 96:26]
  wire [32:0] subRes32 = subed32 - _GEN_0; // @[divR2.scala 96:26]
  wire [31:0] rem32M = subRes32[32] ? subed32[31:0] : subRes32[31:0]; // @[divR2.scala 97:16]
  wire [127:0] div32DividendMux = {64'h0,rem32M,dividendReg[30:0],1'h0}; // @[Cat.scala 29:58]
  wire [64:0] subed64 = dividendReg[127:63]; // @[divR2.scala 91:29]
  wire [64:0] _GEN_1 = {{1'd0}, divisor64Real}; // @[divR2.scala 92:26]
  wire [64:0] subRes64 = subed64 - _GEN_1; // @[divR2.scala 92:26]
  wire [63:0] rem64M = subRes64[64] ? subed64[63:0] : subRes64[63:0]; // @[divR2.scala 93:16]
  wire [127:0] div64DividendMux = {rem64M,dividendReg[62:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_79 = ~subRes32[32]; // @[divR2.scala 104:38]
  wire [63:0] _T_80 = {resReg[62:0],_T_79}; // @[Cat.scala 29:58]
  wire  _T_83 = ~subRes64[64]; // @[divR2.scala 105:38]
  wire [63:0] _T_84 = {resReg[62:0],_T_83}; // @[Cat.scala 29:58]
  wire [63:0] _T_91 = ~resReg; // @[divR2.scala 110:35]
  wire [63:0] _T_93 = _T_91 + 64'h1; // @[divR2.scala 110:53]
  wire [63:0] res64Out = quoSgn64 ? _T_93 : resReg; // @[divR2.scala 110:21]
  wire [63:0] _T_95 = ~dividendReg[127:64]; // @[divR2.scala 111:32]
  wire [63:0] _T_97 = _T_95 + 64'h1; // @[divR2.scala 111:63]
  wire [63:0] rem64Out = _T_1 ? _T_97 : dividendReg[127:64]; // @[divR2.scala 111:20]
  wire [31:0] _T_101 = ~resReg[31:0]; // @[divR2.scala 113:56]
  wire [31:0] _T_103 = _T_101 + 32'h1; // @[divR2.scala 113:79]
  wire [63:0] _T_104 = {32'hffffffff,_T_103}; // @[Cat.scala 29:58]
  wire [63:0] res32out = quoSgn32 ? _T_104 : resReg; // @[divR2.scala 113:21]
  wire [31:0] _T_107 = ~dividendReg[63:32]; // @[divR2.scala 115:56]
  wire [31:0] _T_109 = _T_107 + 32'h1; // @[divR2.scala 115:85]
  wire [63:0] _T_110 = {32'hffffffff,_T_109}; // @[Cat.scala 29:58]
  wire [63:0] _T_113 = {32'h0,dividendReg[63:32]}; // @[Cat.scala 29:58]
  wire [63:0] rem32Out = _T_15 ? _T_110 : _T_113; // @[divR2.scala 115:21]
  assign io_out_valid = stateReg == 2'h3; // @[divR2.scala 123:16]
  assign io_quotient = io_divw ? res32out : res64Out; // @[divR2.scala 119:15]
  assign io_remainder = io_divw ? rem32Out : rem64Out; // @[divR2.scala 120:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {4{`RANDOM}};
  dividendReg = _RAND_2[127:0];
  _RAND_3 = {2{`RANDOM}};
  resReg = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T_42) begin
      if (io_block) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h0;
      end
    end else if (_T_40) begin
      if (_T_37) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h2;
      end
    end else if (_T_38) begin
      if (_T_36) begin
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h1;
      end
    end else if (_T_35) begin
      stateReg <= 2'h2;
    end else if (_T_33) begin
      stateReg <= 2'h1;
    end else begin
      stateReg <= 2'h0;
    end
    if (reset) begin
      cnt <= 6'h0;
    end else if (_T_44) begin
      cnt <= _T_46;
    end else begin
      cnt <= 6'h0;
    end
    if (reset) begin
      dividendReg <= 128'h0;
    end else if (!(_T_42)) begin
      if (_T_40) begin
        dividendReg <= div64DividendMux;
      end else if (_T_38) begin
        dividendReg <= div32DividendMux;
      end else if (_T_35) begin
        dividendReg <= _T_52;
      end else if (_T_33) begin
        dividendReg <= _T_51;
      end else begin
        dividendReg <= 128'h0;
      end
    end
    if (reset) begin
      resReg <= 64'h0;
    end else if (!(_T_42)) begin
      if (_T_40) begin
        resReg <= _T_84;
      end else if (_T_38) begin
        resReg <= _T_80;
      end else begin
        resReg <= 64'h0;
      end
    end
  end
endmodule
module boothSel(
  input  [2:0]   io_y,
  input  [131:0] io_x,
  output [131:0] io_p,
  output         io_c
);
  wire  _T_3 = ~io_y[0]; // @[mul.scala 13:42]
  wire  _T_4 = io_y[1] & _T_3; // @[mul.scala 13:40]
  wire  _T_6 = ~io_y[1]; // @[mul.scala 13:53]
  wire  _T_8 = _T_6 & io_y[0]; // @[mul.scala 13:62]
  wire  _T_9 = _T_4 | _T_8; // @[mul.scala 13:51]
  wire  selNegative = io_y[2] & _T_9; // @[mul.scala 13:29]
  wire  _T_11 = ~io_y[2]; // @[mul.scala 14:21]
  wire  selPositive = _T_11 & _T_9; // @[mul.scala 14:30]
  wire  _T_24 = io_y[2] & _T_6; // @[mul.scala 15:35]
  wire  selDoubleNegative = _T_24 & _T_3; // @[mul.scala 15:46]
  wire  _T_30 = _T_11 & io_y[1]; // @[mul.scala 16:36]
  wire  selDoublePositive = _T_30 & io_y[0]; // @[mul.scala 16:46]
  wire [131:0] _T_33 = selNegative ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _T_34 = ~io_x; // @[mul.scala 18:42]
  wire [131:0] _T_35 = _T_33 & _T_34; // @[mul.scala 18:39]
  wire [131:0] _T_37 = selDoubleNegative ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [130:0] _T_39 = ~io_x[130:0]; // @[mul.scala 19:50]
  wire [131:0] _T_40 = {_T_39,1'h1}; // @[Cat.scala 29:58]
  wire [131:0] _T_41 = _T_37 & _T_40; // @[mul.scala 19:45]
  wire [131:0] _T_42 = _T_35 | _T_41; // @[mul.scala 18:56]
  wire [131:0] _T_44 = selPositive ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _T_45 = _T_44 & io_x; // @[mul.scala 20:39]
  wire [131:0] _T_46 = _T_42 | _T_45; // @[mul.scala 19:79]
  wire [131:0] _T_48 = selDoublePositive ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _T_50 = {io_x[130:0],1'h0}; // @[Cat.scala 29:58]
  wire [131:0] _T_51 = _T_48 & _T_50; // @[mul.scala 21:46]
  assign io_p = _T_46 | _T_51; // @[mul.scala 18:8]
  assign io_c = selDoubleNegative | selNegative; // @[mul.scala 23:8]
endmodule
module add_1(
  input          io_cin,
  input  [131:0] io_a,
  input  [131:0] io_b,
  output [131:0] io_sum
);
  wire [132:0] _T_1 = {1'h0,io_a}; // @[Cat.scala 29:58]
  wire [132:0] _T_2 = {1'h0,io_b}; // @[Cat.scala 29:58]
  wire [132:0] _T_4 = _T_1 + _T_2; // @[add.scala 17:31]
  wire [132:0] _GEN_0 = {{132'd0}, io_cin}; // @[add.scala 17:52]
  wire [132:0] _T_6 = _T_4 + _GEN_0; // @[add.scala 17:52]
  assign io_sum = _T_6[131:0]; // @[add.scala 18:12]
endmodule
module mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [63:0] io_result_low,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] boothIns_io_y; // @[mul.scala 103:24]
  wire [131:0] boothIns_io_x; // @[mul.scala 103:24]
  wire [131:0] boothIns_io_p; // @[mul.scala 103:24]
  wire  boothIns_io_c; // @[mul.scala 103:24]
  wire  addIns_io_cin; // @[mul.scala 105:22]
  wire [131:0] addIns_io_a; // @[mul.scala 105:22]
  wire [131:0] addIns_io_b; // @[mul.scala 105:22]
  wire [131:0] addIns_io_sum; // @[mul.scala 105:22]
  reg [1:0] stateReg; // @[mul.scala 40:25]
  wire  isIdle = stateReg == 2'h0; // @[mul.scala 41:25]
  wire  isMul = stateReg == 2'h1; // @[mul.scala 42:24]
  reg [5:0] cnt; // @[mul.scala 47:20]
  wire  _T = cnt == 6'h20; // @[mul.scala 54:24]
  wire  _T_1 = 2'h0 == stateReg; // @[Mux.scala 80:60]
  wire  _T_3 = 2'h1 == stateReg; // @[Mux.scala 80:60]
  wire  _T_5 = 2'h2 == stateReg; // @[Mux.scala 80:60]
  wire [5:0] _T_8 = cnt + 6'h1; // @[mul.scala 65:25]
  wire [66:0] multiplierEx = {2'h0,io_multiplier,1'h0}; // @[Cat.scala 29:58]
  reg [66:0] multiplierReg; // @[mul.scala 80:30]
  wire  _T_22 = isIdle & io_mul_valid; // @[mul.scala 82:12]
  wire [66:0] _T_24 = {2'h0,multiplierReg[66:2]}; // @[Cat.scala 29:58]
  reg [131:0] multiplicandReg; // @[mul.scala 91:32]
  wire [131:0] _T_28 = {66'h0,2'h0,io_multiplicand}; // @[Cat.scala 29:58]
  wire [131:0] _T_30 = {multiplicandReg[129:0],2'h0}; // @[Cat.scala 29:58]
  reg [131:0] resReg; // @[mul.scala 104:23]
  boothSel boothIns ( // @[mul.scala 103:24]
    .io_y(boothIns_io_y),
    .io_x(boothIns_io_x),
    .io_p(boothIns_io_p),
    .io_c(boothIns_io_c)
  );
  add_1 addIns ( // @[mul.scala 105:22]
    .io_cin(addIns_io_cin),
    .io_a(addIns_io_a),
    .io_b(addIns_io_b),
    .io_sum(addIns_io_sum)
  );
  assign io_out_valid = stateReg == 2'h2; // @[mul.scala 140:16]
  assign io_result_low = resReg[63:0]; // @[mul.scala 137:17]
  assign boothIns_io_y = multiplierReg[2:0]; // @[mul.scala 107:16]
  assign boothIns_io_x = multiplicandReg; // @[mul.scala 108:16]
  assign addIns_io_cin = boothIns_io_c; // @[mul.scala 111:17]
  assign addIns_io_a = boothIns_io_p; // @[mul.scala 110:15]
  assign addIns_io_b = resReg; // @[mul.scala 112:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {3{`RANDOM}};
  multiplierReg = _RAND_2[66:0];
  _RAND_3 = {5{`RANDOM}};
  multiplicandReg = _RAND_3[131:0];
  _RAND_4 = {5{`RANDOM}};
  resReg = _RAND_4[131:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      stateReg <= 2'h0;
    end else if (_T_5) begin
      if (io_block) begin
        stateReg <= 2'h2;
      end else begin
        stateReg <= 2'h0;
      end
    end else if (_T_3) begin
      if (_T) begin
        stateReg <= 2'h2;
      end else begin
        stateReg <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_mul_valid) begin
        stateReg <= 2'h1;
      end else begin
        stateReg <= 2'h0;
      end
    end else begin
      stateReg <= 2'h0;
    end
    if (reset) begin
      cnt <= 6'h0;
    end else if (isMul) begin
      cnt <= _T_8;
    end else begin
      cnt <= 6'h0;
    end
    if (reset) begin
      multiplierReg <= 67'h0;
    end else if (_T_22) begin
      multiplierReg <= multiplierEx;
    end else if (isMul) begin
      multiplierReg <= _T_24;
    end
    if (reset) begin
      multiplicandReg <= 132'h0;
    end else if (_T_22) begin
      multiplicandReg <= _T_28;
    end else if (isMul) begin
      multiplicandReg <= _T_30;
    end
    if (reset) begin
      resReg <= 132'h0;
    end else if (isIdle) begin
      resReg <= 132'h0;
    end else if (isMul) begin
      resReg <= addIns_io_sum;
    end
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_srcA,
  input  [63:0] io_srcB,
  input  [4:0]  io_ALUCtrl,
  output [63:0] io_ALUResult,
  output        block1_0,
  input         block23_0
);
  wire  addIns_io_cin; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_a; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_b; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_sum; // @[ALU.scala 21:22]
  wire  addIns_io_cout; // @[ALU.scala 21:22]
  wire  divR2Ins_clock; // @[ALU.scala 31:23]
  wire  divR2Ins_reset; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_dividend; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_divisor; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_valid; // @[ALU.scala 31:23]
  wire  divR2Ins_io_divw; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_signed; // @[ALU.scala 31:23]
  wire  divR2Ins_io_out_valid; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_quotient; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_remainder; // @[ALU.scala 31:23]
  wire  divR2Ins_io_block; // @[ALU.scala 31:23]
  wire  mulIns_clock; // @[ALU.scala 46:22]
  wire  mulIns_reset; // @[ALU.scala 46:22]
  wire  mulIns_io_mul_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplicand; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplier; // @[ALU.scala 46:22]
  wire  mulIns_io_out_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_result_low; // @[ALU.scala 46:22]
  wire  mulIns_io_block; // @[ALU.scala 46:22]
  wire  _T = io_ALUCtrl == 5'h1; // @[ALU.scala 23:69]
  wire  _T_2 = io_ALUCtrl == 5'h5; // @[ALU.scala 23:69]
  wire  _T_3 = _T | _T_2; // @[ALU.scala 23:56]
  wire  _T_4 = io_ALUCtrl == 5'h10; // @[ALU.scala 23:69]
  wire  _T_5 = _T_3 | _T_4; // @[ALU.scala 23:56]
  wire  _T_7 = _T_5 | _T_2; // @[ALU.scala 23:56]
  wire  _T_8 = io_ALUCtrl == 5'h7; // @[ALU.scala 23:69]
  wire  _T_9 = _T_7 | _T_8; // @[ALU.scala 23:56]
  wire  _T_10 = io_ALUCtrl == 5'h1b; // @[ALU.scala 23:69]
  wire  _T_11 = _T_9 | _T_10; // @[ALU.scala 23:56]
  wire  _T_12 = io_ALUCtrl == 5'h1c; // @[ALU.scala 23:69]
  wire  sub = _T_11 | _T_12; // @[ALU.scala 23:56]
  wire [63:0] srcBInv = ~io_srcB; // @[ALU.scala 24:18]
  wire  _T_14 = io_ALUCtrl == 5'h11; // @[ALU.scala 33:79]
  wire  _T_16 = io_ALUCtrl == 5'h12; // @[ALU.scala 33:79]
  wire  _T_17 = _T_14 | _T_16; // @[ALU.scala 33:66]
  wire  _T_18 = io_ALUCtrl == 5'h14; // @[ALU.scala 33:79]
  wire  _T_19 = _T_17 | _T_18; // @[ALU.scala 33:66]
  wire  _T_20 = io_ALUCtrl == 5'h15; // @[ALU.scala 33:79]
  wire  _T_21 = _T_19 | _T_20; // @[ALU.scala 33:66]
  wire  _T_22 = io_ALUCtrl == 5'h17; // @[ALU.scala 33:79]
  wire  _T_23 = _T_21 | _T_22; // @[ALU.scala 33:66]
  wire  _T_24 = io_ALUCtrl == 5'h18; // @[ALU.scala 33:79]
  wire  _T_25 = _T_23 | _T_24; // @[ALU.scala 33:66]
  wire  _T_26 = io_ALUCtrl == 5'h19; // @[ALU.scala 33:79]
  wire  _T_27 = _T_25 | _T_26; // @[ALU.scala 33:66]
  wire  _T_28 = io_ALUCtrl == 5'h1d; // @[ALU.scala 33:79]
  wire  _T_39 = _T_18 | _T_20; // @[ALU.scala 37:68]
  wire  _T_41 = _T_39 | _T_24; // @[ALU.scala 37:68]
  wire [63:0] srcAUSignW = {32'h0,io_srcA[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] srcBUSignW = {32'h0,io_srcB[31:0]}; // @[Cat.scala 29:58]
  wire  _T_45 = io_ALUCtrl == 5'h13; // @[ALU.scala 50:79]
  wire  _T_47 = io_ALUCtrl == 5'h16; // @[ALU.scala 50:79]
  wire [5:0] shamt = io_srcB[5:0]; // @[ALU.scala 61:22]
  wire [63:0] _T_53 = $signed(io_srcA) >>> shamt; // @[ALU.scala 65:42]
  wire [63:0] _T_54 = io_srcA >> shamt; // @[ALU.scala 66:25]
  wire [126:0] _GEN_0 = {{63'd0}, io_srcA}; // @[ALU.scala 67:25]
  wire [126:0] _T_55 = _GEN_0 << shamt; // @[ALU.scala 67:25]
  wire  _T_57 = ~addIns_io_cout; // @[ALU.scala 69:16]
  wire [63:0] _T_58 = io_srcA & io_srcB; // @[ALU.scala 70:25]
  wire [63:0] _T_59 = io_srcA | io_srcB; // @[ALU.scala 71:24]
  wire [63:0] _T_60 = io_srcA ^ io_srcB; // @[ALU.scala 72:25]
  wire  _T_61 = io_srcA != io_srcB; // @[ALU.scala 73:32]
  wire [63:0] _T_62 = {63'h0,_T_61}; // @[Cat.scala 29:58]
  wire [31:0] _T_64 = io_srcA[31:0] >> shamt; // @[ALU.scala 74:48]
  wire [31:0] _T_67 = _T_64[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_68 = {_T_67,_T_64}; // @[Cat.scala 29:58]
  wire [31:0] _T_72 = addIns_io_sum[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_73 = {_T_72,addIns_io_sum[31:0]}; // @[Cat.scala 29:58]
  wire [94:0] _GEN_1 = {{63'd0}, io_srcA[31:0]}; // @[ALU.scala 76:48]
  wire [94:0] _T_75 = _GEN_1 << shamt; // @[ALU.scala 76:48]
  wire [31:0] _T_79 = _T_75[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_80 = {_T_79,_T_75[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_82 = io_srcA[31:0]; // @[ALU.scala 77:41]
  wire [31:0] _T_84 = $signed(_T_82) >>> shamt; // @[ALU.scala 77:65]
  wire [31:0] _T_87 = _T_84[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_88 = {_T_87,_T_84}; // @[Cat.scala 29:58]
  wire [31:0] _T_97 = divR2Ins_io_quotient[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_98 = {_T_97,divR2Ins_io_quotient[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_102 = divR2Ins_io_remainder[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_103 = {_T_102,divR2Ins_io_remainder[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_107 = mulIns_io_result_low[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_108 = {_T_107,mulIns_io_result_low[31:0]}; // @[Cat.scala 29:58]
  wire  _T_119 = io_srcA == io_srcB; // @[ALU.scala 88:24]
  wire  _T_121 = ~addIns_io_sum[63]; // @[ALU.scala 91:16]
  wire  _T_122 = 5'h0 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_123 = _T_122 ? addIns_io_sum : 64'h0; // @[Mux.scala 80:57]
  wire  _T_124 = 5'h1 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_125 = _T_124 ? addIns_io_sum : _T_123; // @[Mux.scala 80:57]
  wire  _T_126 = 5'h9 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_127 = _T_126 ? _T_53 : _T_125; // @[Mux.scala 80:57]
  wire  _T_128 = 5'h8 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [63:0] _T_129 = _T_128 ? _T_54 : _T_127; // @[Mux.scala 80:57]
  wire  _T_130 = 5'h6 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_131 = _T_130 ? _T_55 : {{63'd0}, _T_129}; // @[Mux.scala 80:57]
  wire  _T_132 = 5'h5 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_133 = _T_132 ? {{126'd0}, addIns_io_sum[63]} : _T_131; // @[Mux.scala 80:57]
  wire  _T_134 = 5'h7 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_135 = _T_134 ? {{126'd0}, _T_57} : _T_133; // @[Mux.scala 80:57]
  wire  _T_136 = 5'h2 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_137 = _T_136 ? {{63'd0}, _T_58} : _T_135; // @[Mux.scala 80:57]
  wire  _T_138 = 5'h3 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_139 = _T_138 ? {{63'd0}, _T_59} : _T_137; // @[Mux.scala 80:57]
  wire  _T_140 = 5'h4 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_141 = _T_140 ? {{63'd0}, _T_60} : _T_139; // @[Mux.scala 80:57]
  wire  _T_142 = 5'hb == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_143 = _T_142 ? {{63'd0}, _T_62} : _T_141; // @[Mux.scala 80:57]
  wire  _T_144 = 5'hc == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_145 = _T_144 ? {{63'd0}, _T_68} : _T_143; // @[Mux.scala 80:57]
  wire  _T_146 = 5'hd == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_147 = _T_146 ? {{63'd0}, _T_73} : _T_145; // @[Mux.scala 80:57]
  wire  _T_148 = 5'he == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_149 = _T_148 ? {{63'd0}, _T_80} : _T_147; // @[Mux.scala 80:57]
  wire  _T_150 = 5'hf == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_151 = _T_150 ? {{63'd0}, _T_88} : _T_149; // @[Mux.scala 80:57]
  wire  _T_152 = 5'h10 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_153 = _T_152 ? {{63'd0}, _T_73} : _T_151; // @[Mux.scala 80:57]
  wire  _T_154 = 5'h11 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_155 = _T_154 ? {{63'd0}, _T_98} : _T_153; // @[Mux.scala 80:57]
  wire  _T_156 = 5'h12 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_157 = _T_156 ? {{63'd0}, _T_103} : _T_155; // @[Mux.scala 80:57]
  wire  _T_158 = 5'h13 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_159 = _T_158 ? {{63'd0}, _T_108} : _T_157; // @[Mux.scala 80:57]
  wire  _T_160 = 5'h14 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_161 = _T_160 ? {{63'd0}, _T_103} : _T_159; // @[Mux.scala 80:57]
  wire  _T_162 = 5'h15 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_163 = _T_162 ? {{63'd0}, _T_98} : _T_161; // @[Mux.scala 80:57]
  wire  _T_164 = 5'h16 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_165 = _T_164 ? {{63'd0}, mulIns_io_result_low} : _T_163; // @[Mux.scala 80:57]
  wire  _T_166 = 5'h17 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_167 = _T_166 ? {{63'd0}, divR2Ins_io_quotient} : _T_165; // @[Mux.scala 80:57]
  wire  _T_168 = 5'h18 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_169 = _T_168 ? {{63'd0}, divR2Ins_io_remainder} : _T_167; // @[Mux.scala 80:57]
  wire  _T_170 = 5'h19 == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_171 = _T_170 ? {{63'd0}, divR2Ins_io_quotient} : _T_169; // @[Mux.scala 80:57]
  wire  _T_172 = 5'h1a == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_173 = _T_172 ? {{126'd0}, _T_119} : _T_171; // @[Mux.scala 80:57]
  wire  _T_174 = 5'h1b == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_175 = _T_174 ? {{126'd0}, addIns_io_cout} : _T_173; // @[Mux.scala 80:57]
  wire  _T_176 = 5'h1c == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_177 = _T_176 ? {{126'd0}, _T_121} : _T_175; // @[Mux.scala 80:57]
  wire  _T_178 = 5'h1d == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_179 = _T_178 ? {{63'd0}, divR2Ins_io_remainder} : _T_177; // @[Mux.scala 80:57]
  wire  _T_180 = 5'ha == io_ALUCtrl; // @[Mux.scala 80:60]
  wire [126:0] _T_181 = _T_180 ? {{63'd0}, io_srcA} : _T_179; // @[Mux.scala 80:57]
  wire  _T_182 = ~divR2Ins_io_out_valid; // @[ALU.scala 98:38]
  wire  _T_183 = divR2Ins_io_div_valid & _T_182; // @[ALU.scala 98:35]
  wire  _T_184 = ~mulIns_io_out_valid; // @[ALU.scala 98:87]
  wire  _T_185 = mulIns_io_mul_valid & _T_184; // @[ALU.scala 98:84]
  wire  _T_186 = _T_183 | _T_185; // @[ALU.scala 98:61]
  wire  block1 = _T_186; // @[ALU.scala 97:20 ALU.scala 98:10]
  add addIns ( // @[ALU.scala 21:22]
    .io_cin(addIns_io_cin),
    .io_a(addIns_io_a),
    .io_b(addIns_io_b),
    .io_sum(addIns_io_sum),
    .io_cout(addIns_io_cout)
  );
  divR2 divR2Ins ( // @[ALU.scala 31:23]
    .clock(divR2Ins_clock),
    .reset(divR2Ins_reset),
    .io_dividend(divR2Ins_io_dividend),
    .io_divisor(divR2Ins_io_divisor),
    .io_div_valid(divR2Ins_io_div_valid),
    .io_divw(divR2Ins_io_divw),
    .io_div_signed(divR2Ins_io_div_signed),
    .io_out_valid(divR2Ins_io_out_valid),
    .io_quotient(divR2Ins_io_quotient),
    .io_remainder(divR2Ins_io_remainder),
    .io_block(divR2Ins_io_block)
  );
  mul mulIns ( // @[ALU.scala 46:22]
    .clock(mulIns_clock),
    .reset(mulIns_reset),
    .io_mul_valid(mulIns_io_mul_valid),
    .io_multiplicand(mulIns_io_multiplicand),
    .io_multiplier(mulIns_io_multiplier),
    .io_out_valid(mulIns_io_out_valid),
    .io_result_low(mulIns_io_result_low),
    .io_block(mulIns_io_block)
  );
  assign io_ALUResult = _T_181[63:0]; // @[ALU.scala 95:16]
  assign block1_0 = block1;
  assign addIns_io_cin = _T_11 | _T_12; // @[ALU.scala 25:17]
  assign addIns_io_a = io_srcA; // @[ALU.scala 26:15]
  assign addIns_io_b = sub ? srcBInv : io_srcB; // @[ALU.scala 28:15]
  assign divR2Ins_clock = clock;
  assign divR2Ins_reset = reset;
  assign divR2Ins_io_dividend = io_srcA; // @[ALU.scala 38:24]
  assign divR2Ins_io_divisor = io_srcB; // @[ALU.scala 39:23]
  assign divR2Ins_io_div_valid = _T_27 | _T_28; // @[ALU.scala 40:25]
  assign divR2Ins_io_divw = _T_19 | _T_20; // @[ALU.scala 41:20]
  assign divR2Ins_io_div_signed = _T_41 | _T_26; // @[ALU.scala 42:26]
  assign divR2Ins_io_block = block23_0; // @[ALU.scala 111:21]
  assign mulIns_clock = clock;
  assign mulIns_reset = reset;
  assign mulIns_io_mul_valid = _T_45 | _T_47; // @[ALU.scala 55:23]
  assign mulIns_io_multiplicand = _T_45 ? srcAUSignW : io_srcA; // @[ALU.scala 56:26]
  assign mulIns_io_multiplier = _T_45 ? srcBUSignW : io_srcB; // @[ALU.scala 57:24]
  assign mulIns_io_block = block23_0; // @[ALU.scala 110:19]
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_csrrwen,
  input         io_csrswen,
  input         io_csrrsien,
  input         io_csrrcien,
  input         io_csrrcen,
  input         io_csrrwien,
  input         io_ecall,
  input  [63:0] io_rs1,
  input  [11:0] io_imme,
  input  [63:0] io_pc,
  input  [4:0]  io_uimm,
  output [63:0] io_rd,
  output [63:0] io_mtvec,
  output [63:0] io_mepc,
  input         io_mret,
  input         intrTimeCnt_0,
  output        startTimeCnt_0,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_pc != 64'h0; // @[CSR.scala 37:35]
  wire  intr = intrTimeCnt_0 & _T; // @[CSR.scala 37:26]
  wire  _T_1 = io_csrrwen | io_csrswen; // @[CSR.scala 51:26]
  wire  _T_2 = _T_1 | io_csrrcen; // @[CSR.scala 51:38]
  wire  _T_3 = _T_2 | io_csrrsien; // @[CSR.scala 51:52]
  wire  _T_4 = _T_3 | io_csrrcien; // @[CSR.scala 51:67]
  wire  csren = _T_4 | io_csrrwien; // @[CSR.scala 51:82]
  wire [5:0] sel1H = {io_csrrwien,io_csrrcien,io_csrrsien,io_csrrcen,io_csrswen,io_csrrwen}; // @[Cat.scala 29:58]
  wire [63:0] uimmext = {59'h0,io_uimm}; // @[Cat.scala 29:58]
  wire  _T_9 = io_imme == 12'h341; // @[CSR.scala 55:48]
  wire  _T_10 = csren & _T_9; // @[CSR.scala 55:36]
  wire  _T_11 = io_ecall | _T_10; // @[CSR.scala 55:25]
  wire  mepcen = _T_11 | intr; // @[CSR.scala 55:58]
  wire  _T_12 = io_ecall | intr; // @[CSR.scala 58:14]
  reg [63:0] mepcins; // @[Reg.scala 27:20]
  wire [63:0] _T_13 = io_rs1 | mepcins; // @[CSR.scala 64:15]
  wire [63:0] _T_14 = ~io_rs1; // @[CSR.scala 65:10]
  wire [63:0] _T_15 = _T_14 & mepcins; // @[CSR.scala 65:28]
  wire [63:0] _T_16 = uimmext | mepcins; // @[CSR.scala 66:17]
  wire [63:0] _T_17 = ~uimmext; // @[CSR.scala 67:10]
  wire [63:0] _T_18 = _T_17 & mepcins; // @[CSR.scala 67:29]
  wire [63:0] _T_25 = sel1H[0] ? io_rs1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_26 = sel1H[1] ? _T_13 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_27 = sel1H[2] ? _T_15 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_28 = sel1H[3] ? _T_16 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_29 = sel1H[4] ? _T_18 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_30 = sel1H[5] ? uimmext : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_31 = _T_25 | _T_26; // @[Mux.scala 27:72]
  wire [63:0] _T_32 = _T_31 | _T_27; // @[Mux.scala 27:72]
  wire [63:0] _T_33 = _T_32 | _T_28; // @[Mux.scala 27:72]
  wire [63:0] _T_34 = _T_33 | _T_29; // @[Mux.scala 27:72]
  wire [63:0] _T_35 = _T_34 | _T_30; // @[Mux.scala 27:72]
  wire  _T_37 = block1_0 | block23_0; // @[CSR.scala 72:56]
  wire  _T_38 = ~_T_37; // @[CSR.scala 72:47]
  wire  _T_39 = mepcen & _T_38; // @[CSR.scala 72:44]
  wire  _T_41 = io_imme == 12'h342; // @[CSR.scala 74:49]
  wire  _T_42 = csren & _T_41; // @[CSR.scala 74:37]
  wire  _T_43 = io_ecall | _T_42; // @[CSR.scala 74:27]
  wire  mcauseen = _T_43 | intr; // @[CSR.scala 74:61]
  reg [63:0] mcauseins; // @[Reg.scala 27:20]
  wire [63:0] _T_44 = io_rs1 | mcauseins; // @[CSR.scala 86:16]
  wire [63:0] _T_46 = _T_14 & mcauseins; // @[CSR.scala 87:28]
  wire [63:0] _T_47 = uimmext | mcauseins; // @[CSR.scala 88:17]
  wire [63:0] _T_49 = _T_17 & mcauseins; // @[CSR.scala 89:29]
  wire [63:0] _T_57 = sel1H[1] ? _T_44 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_58 = sel1H[2] ? _T_46 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_59 = sel1H[3] ? _T_47 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_60 = sel1H[4] ? _T_49 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_62 = _T_25 | _T_57; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_62 | _T_58; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = _T_63 | _T_59; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = _T_64 | _T_60; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = _T_65 | _T_30; // @[Mux.scala 27:72]
  wire  _T_71 = mcauseen & _T_38; // @[CSR.scala 94:50]
  wire  _T_73 = io_imme == 12'h305; // @[CSR.scala 96:37]
  wire  mtvecen = csren & _T_73; // @[CSR.scala 96:25]
  reg [63:0] mtvecins; // @[Reg.scala 27:20]
  wire [63:0] _T_74 = io_rs1 | mtvecins; // @[CSR.scala 102:14]
  wire [63:0] _T_76 = _T_14 & mtvecins; // @[CSR.scala 103:26]
  wire [63:0] _T_77 = uimmext | mtvecins; // @[CSR.scala 104:15]
  wire [63:0] _T_79 = _T_17 & mtvecins; // @[CSR.scala 105:27]
  wire [63:0] _T_87 = sel1H[1] ? _T_74 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_88 = sel1H[2] ? _T_76 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_89 = sel1H[3] ? _T_77 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_90 = sel1H[4] ? _T_79 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_92 = _T_25 | _T_87; // @[Mux.scala 27:72]
  wire [63:0] _T_93 = _T_92 | _T_88; // @[Mux.scala 27:72]
  wire [63:0] _T_94 = _T_93 | _T_89; // @[Mux.scala 27:72]
  wire [63:0] _T_95 = _T_94 | _T_90; // @[Mux.scala 27:72]
  wire [63:0] mtvecval = _T_95 | _T_30; // @[Mux.scala 27:72]
  wire  _T_98 = _T_37 | intr; // @[CSR.scala 109:70]
  wire  _T_99 = ~_T_98; // @[CSR.scala 109:50]
  wire  _T_100 = mtvecen & _T_99; // @[CSR.scala 109:47]
  wire  _T_102 = io_imme == 12'h300; // @[CSR.scala 111:40]
  wire  _T_103 = csren & _T_102; // @[CSR.scala 111:28]
  wire  _T_104 = _T_103 | io_ecall; // @[CSR.scala 111:54]
  wire  _T_105 = _T_104 | intr; // @[CSR.scala 111:65]
  wire  mstatusen = _T_105 | io_mret; // @[CSR.scala 111:73]
  reg [63:0] mstatusins; // @[Reg.scala 27:20]
  wire [63:0] _T_114 = {mstatusins[63:8],mstatusins[3],mstatusins[6:4],1'h0,mstatusins[2:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_122 = {mstatusins[63:8],1'h1,mstatusins[6:4],mstatusins[7],mstatusins[2:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_123 = io_rs1 | mstatusins; // @[CSR.scala 124:14]
  wire [63:0] _T_125 = _T_14 & mstatusins; // @[CSR.scala 125:26]
  wire [63:0] _T_126 = uimmext | mstatusins; // @[CSR.scala 126:15]
  wire [63:0] _T_128 = _T_17 & mstatusins; // @[CSR.scala 127:27]
  wire [63:0] _T_136 = sel1H[1] ? _T_123 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_137 = sel1H[2] ? _T_125 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_138 = sel1H[3] ? _T_126 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_139 = sel1H[4] ? _T_128 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_141 = _T_25 | _T_136; // @[Mux.scala 27:72]
  wire [63:0] _T_142 = _T_141 | _T_137; // @[Mux.scala 27:72]
  wire [63:0] _T_143 = _T_142 | _T_138; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_143 | _T_139; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_144 | _T_30; // @[Mux.scala 27:72]
  wire  _T_150 = mstatusen & _T_38; // @[CSR.scala 148:73]
  wire  _T_152 = io_imme == 12'h304; // @[CSR.scala 150:36]
  wire  miecen = csren & _T_152; // @[CSR.scala 150:24]
  reg [63:0] mieins; // @[Reg.scala 27:20]
  wire [63:0] _T_153 = io_rs1 | mieins; // @[CSR.scala 156:14]
  wire [63:0] _T_155 = _T_14 & mieins; // @[CSR.scala 157:26]
  wire [63:0] _T_156 = uimmext | mieins; // @[CSR.scala 158:15]
  wire [63:0] _T_158 = _T_17 & mieins; // @[CSR.scala 159:27]
  wire [63:0] _T_166 = sel1H[1] ? _T_153 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_167 = sel1H[2] ? _T_155 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_168 = sel1H[3] ? _T_156 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_169 = sel1H[4] ? _T_158 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_171 = _T_25 | _T_166; // @[Mux.scala 27:72]
  wire [63:0] _T_172 = _T_171 | _T_167; // @[Mux.scala 27:72]
  wire [63:0] _T_173 = _T_172 | _T_168; // @[Mux.scala 27:72]
  wire [63:0] _T_174 = _T_173 | _T_169; // @[Mux.scala 27:72]
  wire [63:0] mieval = _T_174 | _T_30; // @[Mux.scala 27:72]
  wire  _T_179 = miecen & _T_99; // @[CSR.scala 163:41]
  wire  _T_181 = io_imme == 12'h344; // @[CSR.scala 165:35]
  wire  _T_182 = csren & _T_181; // @[CSR.scala 165:23]
  wire  mipcen = _T_182 | intr; // @[CSR.scala 165:45]
  reg [63:0] mipins; // @[Reg.scala 27:20]
  wire [63:0] _T_186 = {mipins[63:8],1'h1,mipins[6:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_187 = io_rs1 | mipins; // @[CSR.scala 174:14]
  wire [63:0] _T_189 = _T_14 & mipins; // @[CSR.scala 175:26]
  wire [63:0] _T_190 = uimmext | mipins; // @[CSR.scala 176:15]
  wire [63:0] _T_192 = _T_17 & mipins; // @[CSR.scala 177:27]
  wire [63:0] _T_200 = sel1H[1] ? _T_187 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_201 = sel1H[2] ? _T_189 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_202 = sel1H[3] ? _T_190 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_203 = sel1H[4] ? _T_192 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_205 = _T_25 | _T_200; // @[Mux.scala 27:72]
  wire [63:0] _T_206 = _T_205 | _T_201; // @[Mux.scala 27:72]
  wire [63:0] _T_207 = _T_206 | _T_202; // @[Mux.scala 27:72]
  wire [63:0] _T_208 = _T_207 | _T_203; // @[Mux.scala 27:72]
  wire [63:0] _T_209 = _T_208 | _T_30; // @[Mux.scala 27:72]
  wire  _T_213 = mipcen & _T_38; // @[CSR.scala 181:42]
  wire  _T_215 = 12'h341 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_216 = _T_215 ? mepcins : 64'h0; // @[Mux.scala 80:57]
  wire  _T_217 = 12'h342 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_218 = _T_217 ? mcauseins : _T_216; // @[Mux.scala 80:57]
  wire  _T_219 = 12'h305 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_220 = _T_219 ? mtvecins : _T_218; // @[Mux.scala 80:57]
  wire  _T_221 = 12'h300 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_222 = _T_221 ? mstatusins : _T_220; // @[Mux.scala 80:57]
  wire  _T_223 = 12'h304 == io_imme; // @[Mux.scala 80:60]
  wire [63:0] _T_224 = _T_223 ? mieins : _T_222; // @[Mux.scala 80:57]
  wire  _T_225 = 12'h344 == io_imme; // @[Mux.scala 80:60]
  wire  _T_229 = mieins[7] & mstatusins[3]; // @[CSR.scala 239:29]
  wire  startTimeCnt = _T_229; // @[CSR.scala 238:26 CSR.scala 239:16]
  assign io_rd = _T_225 ? mipins : _T_224; // @[CSR.scala 219:9]
  assign io_mtvec = mtvecins; // @[CSR.scala 235:12]
  assign io_mepc = mepcins; // @[CSR.scala 236:11]
  assign startTimeCnt_0 = startTimeCnt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mepcins = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcauseins = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvecins = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatusins = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mieins = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mipins = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mepcins <= 64'h0;
    end else if (_T_39) begin
      if (_T_12) begin
        mepcins <= io_pc;
      end else begin
        mepcins <= _T_35;
      end
    end
    if (reset) begin
      mcauseins <= 64'h0;
    end else if (_T_71) begin
      if (intr) begin
        mcauseins <= 64'h8000000000000007;
      end else if (io_ecall) begin
        mcauseins <= 64'hb;
      end else begin
        mcauseins <= _T_66;
      end
    end
    if (reset) begin
      mtvecins <= 64'h0;
    end else if (_T_100) begin
      mtvecins <= mtvecval;
    end
    if (reset) begin
      mstatusins <= 64'ha00001800;
    end else if (_T_150) begin
      if (_T_12) begin
        mstatusins <= _T_114;
      end else if (io_mret) begin
        mstatusins <= _T_122;
      end else begin
        mstatusins <= _T_145;
      end
    end
    if (reset) begin
      mieins <= 64'h0;
    end else if (_T_179) begin
      mieins <= mieval;
    end
    if (reset) begin
      mipins <= 64'h0;
    end else if (_T_213) begin
      if (intr) begin
        mipins <= _T_186;
      end else begin
        mipins <= _T_209;
      end
    end
  end
endmodule
module dnpcGen(
  input         io_npcSrc,
  input  [31:0] io_pc,
  input  [31:0] io_imme,
  input  [31:0] io_rd,
  output [31:0] io_dnpc
);
  wire  _T = ~io_npcSrc; // @[dnpcGen.scala 15:28]
  wire [31:0] src1 = _T ? io_rd : io_pc; // @[dnpcGen.scala 15:17]
  assign io_dnpc = io_imme + src1; // @[dnpcGen.scala 16:11]
endmodule
module memData(
  input  [63:0] io_rdata,
  output [63:0] io_rdata_ext,
  input  [2:0]  io_memReadNum
);
  wire [55:0] _T_3 = io_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_4 = {_T_3,io_rdata[7:0]}; // @[Cat.scala 29:58]
  wire [47:0] _T_8 = io_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_9 = {_T_8,io_rdata[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_13 = io_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_14 = {_T_13,io_rdata[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_16 = {56'h0,io_rdata[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_18 = {48'h0,io_rdata[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_20 = {32'h0,io_rdata[31:0]}; // @[Cat.scala 29:58]
  wire  _T_21 = 3'h0 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_22 = _T_21 ? _T_4 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_23 = 3'h1 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_24 = _T_23 ? _T_9 : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 3'h2 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_26 = _T_25 ? _T_14 : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 3'h3 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_28 = _T_27 ? io_rdata : _T_26; // @[Mux.scala 80:57]
  wire  _T_29 = 3'h4 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_30 = _T_29 ? _T_16 : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 3'h5 == io_memReadNum; // @[Mux.scala 80:60]
  wire [63:0] _T_32 = _T_31 ? _T_18 : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 3'h6 == io_memReadNum; // @[Mux.scala 80:60]
  assign io_rdata_ext = _T_33 ? _T_20 : _T_32; // @[memData.scala 13:16]
endmodule
module execute(
  input         clock,
  input         reset,
  input  [1:0]  io_AluSrc1,
  input  [1:0]  io_AluSrc2,
  input  [4:0]  io_ALUCtrl,
  input         io_dnpcSrc,
  input  [1:0]  io_ResultSrc,
  input  [2:0]  io_memReadNum,
  input  [63:0] io_dataId_imme,
  input  [63:0] io_dataId_dOut1,
  input  [63:0] io_dataId_dOut2,
  output [63:0] io_dataId_dIn,
  output [63:0] io_dataOut_ALUResOut,
  output [63:0] io_dataOut_wdata,
  input  [63:0] io_dataOut_rdata,
  output        io_brTake,
  input  [31:0] io_pc,
  input  [31:0] io_snpc,
  output [31:0] io_dnpc,
  input         io_CSRCtrlIf_csrrwen,
  input         io_CSRCtrlIf_csrswen,
  input         io_CSRCtrlIf_csrrsien,
  input         io_CSRCtrlIf_csrrcien,
  input         io_CSRCtrlIf_csrrcen,
  input         io_CSRCtrlIf_csrrwien,
  input         io_CSRCtrlIf_ecall,
  input         io_CSRCtrlIf_rfen,
  input         io_CSRCtrlIf_mepc2pc,
  input  [4:0]  io_uimm,
  input  [63:0] io_aluResIn,
  input  [1:0]  io_forwardA,
  input  [1:0]  io_forwardB,
  input  [63:0] io_aluRes1,
  input  [63:0] io_aluRes3,
  input         intrTimeCnt_0,
  output        startTimeCnt,
  output        block1,
  input         block23
);
  wire  ALU_clock; // @[execute.scala 96:19]
  wire  ALU_reset; // @[execute.scala 96:19]
  wire [63:0] ALU_io_srcA; // @[execute.scala 96:19]
  wire [63:0] ALU_io_srcB; // @[execute.scala 96:19]
  wire [4:0] ALU_io_ALUCtrl; // @[execute.scala 96:19]
  wire [63:0] ALU_io_ALUResult; // @[execute.scala 96:19]
  wire  ALU_block1_0; // @[execute.scala 96:19]
  wire  ALU_block23_0; // @[execute.scala 96:19]
  wire  csr_ins_clock; // @[execute.scala 103:23]
  wire  csr_ins_reset; // @[execute.scala 103:23]
  wire  csr_ins_io_csrrwen; // @[execute.scala 103:23]
  wire  csr_ins_io_csrswen; // @[execute.scala 103:23]
  wire  csr_ins_io_csrrsien; // @[execute.scala 103:23]
  wire  csr_ins_io_csrrcien; // @[execute.scala 103:23]
  wire  csr_ins_io_csrrcen; // @[execute.scala 103:23]
  wire  csr_ins_io_csrrwien; // @[execute.scala 103:23]
  wire  csr_ins_io_ecall; // @[execute.scala 103:23]
  wire [63:0] csr_ins_io_rs1; // @[execute.scala 103:23]
  wire [11:0] csr_ins_io_imme; // @[execute.scala 103:23]
  wire [63:0] csr_ins_io_pc; // @[execute.scala 103:23]
  wire [4:0] csr_ins_io_uimm; // @[execute.scala 103:23]
  wire [63:0] csr_ins_io_rd; // @[execute.scala 103:23]
  wire [63:0] csr_ins_io_mtvec; // @[execute.scala 103:23]
  wire [63:0] csr_ins_io_mepc; // @[execute.scala 103:23]
  wire  csr_ins_io_mret; // @[execute.scala 103:23]
  wire  csr_ins_intrTimeCnt_0; // @[execute.scala 103:23]
  wire  csr_ins_startTimeCnt_0; // @[execute.scala 103:23]
  wire  csr_ins_block1_0; // @[execute.scala 103:23]
  wire  csr_ins_block23_0; // @[execute.scala 103:23]
  wire  dnpcGenIns_io_npcSrc; // @[execute.scala 123:26]
  wire [31:0] dnpcGenIns_io_pc; // @[execute.scala 123:26]
  wire [31:0] dnpcGenIns_io_imme; // @[execute.scala 123:26]
  wire [31:0] dnpcGenIns_io_rd; // @[execute.scala 123:26]
  wire [31:0] dnpcGenIns_io_dnpc; // @[execute.scala 123:26]
  wire [63:0] memData_ins_io_rdata; // @[execute.scala 148:27]
  wire [63:0] memData_ins_io_rdata_ext; // @[execute.scala 148:27]
  wire [2:0] memData_ins_io_memReadNum; // @[execute.scala 148:27]
  wire  _T = 2'h2 == io_forwardA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? io_aluRes1 : io_dataId_dOut1; // @[Mux.scala 80:57]
  wire  _T_2 = 2'h1 == io_forwardA; // @[Mux.scala 80:60]
  wire  _T_30 = 2'h2 == io_ResultSrc; // @[Mux.scala 80:60]
  wire  _T_28 = 2'h1 == io_ResultSrc; // @[Mux.scala 80:60]
  wire [63:0] _T_29 = _T_28 ? {{32'd0}, io_snpc} : io_aluResIn; // @[Mux.scala 80:57]
  wire [63:0] dinMux = _T_30 ? memData_ins_io_rdata_ext : _T_29; // @[Mux.scala 80:57]
  wire [63:0] _T_3 = _T_2 ? dinMux : _T_1; // @[Mux.scala 80:57]
  wire  _T_4 = 2'h3 == io_forwardA; // @[Mux.scala 80:60]
  wire [63:0] dOut1 = _T_4 ? io_aluRes3 : _T_3; // @[Mux.scala 80:57]
  wire  _T_5 = 2'h0 == io_AluSrc1; // @[Mux.scala 80:60]
  wire [63:0] _T_6 = _T_5 ? dOut1 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_7 = 2'h1 == io_AluSrc1; // @[Mux.scala 80:60]
  wire [63:0] _T_8 = _T_7 ? io_dataId_imme : _T_6; // @[Mux.scala 80:57]
  wire  _T_9 = 2'h2 == io_AluSrc1; // @[Mux.scala 80:60]
  wire  _T_10 = 2'h2 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] _T_11 = _T_10 ? io_aluRes1 : io_dataId_dOut2; // @[Mux.scala 80:57]
  wire  _T_12 = 2'h1 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] _T_13 = _T_12 ? dinMux : _T_11; // @[Mux.scala 80:57]
  wire  _T_14 = 2'h3 == io_forwardB; // @[Mux.scala 80:60]
  wire [63:0] dOut2 = _T_14 ? io_aluRes3 : _T_13; // @[Mux.scala 80:57]
  wire  _T_15 = 2'h0 == io_AluSrc2; // @[Mux.scala 80:60]
  wire [63:0] _T_16 = _T_15 ? dOut2 : 64'h0; // @[Mux.scala 80:57]
  wire  _T_17 = 2'h1 == io_AluSrc2; // @[Mux.scala 80:60]
  wire [63:0] _T_18 = _T_17 ? io_dataId_imme : _T_16; // @[Mux.scala 80:57]
  wire  _T_19 = 2'h2 == io_AluSrc2; // @[Mux.scala 80:60]
  wire  _T_21 = io_CSRCtrlIf_ecall | intrTimeCnt_0; // @[execute.scala 134:37]
  wire [63:0] _T_22 = io_CSRCtrlIf_mepc2pc ? csr_ins_io_mepc : {{32'd0}, dnpcGenIns_io_dnpc}; // @[execute.scala 134:72]
  wire [63:0] _T_23 = _T_21 ? csr_ins_io_mtvec : _T_22; // @[execute.scala 134:17]
  ALU ALU ( // @[execute.scala 96:19]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_srcA(ALU_io_srcA),
    .io_srcB(ALU_io_srcB),
    .io_ALUCtrl(ALU_io_ALUCtrl),
    .io_ALUResult(ALU_io_ALUResult),
    .block1_0(ALU_block1_0),
    .block23_0(ALU_block23_0)
  );
  CSR csr_ins ( // @[execute.scala 103:23]
    .clock(csr_ins_clock),
    .reset(csr_ins_reset),
    .io_csrrwen(csr_ins_io_csrrwen),
    .io_csrswen(csr_ins_io_csrswen),
    .io_csrrsien(csr_ins_io_csrrsien),
    .io_csrrcien(csr_ins_io_csrrcien),
    .io_csrrcen(csr_ins_io_csrrcen),
    .io_csrrwien(csr_ins_io_csrrwien),
    .io_ecall(csr_ins_io_ecall),
    .io_rs1(csr_ins_io_rs1),
    .io_imme(csr_ins_io_imme),
    .io_pc(csr_ins_io_pc),
    .io_uimm(csr_ins_io_uimm),
    .io_rd(csr_ins_io_rd),
    .io_mtvec(csr_ins_io_mtvec),
    .io_mepc(csr_ins_io_mepc),
    .io_mret(csr_ins_io_mret),
    .intrTimeCnt_0(csr_ins_intrTimeCnt_0),
    .startTimeCnt_0(csr_ins_startTimeCnt_0),
    .block1_0(csr_ins_block1_0),
    .block23_0(csr_ins_block23_0)
  );
  dnpcGen dnpcGenIns ( // @[execute.scala 123:26]
    .io_npcSrc(dnpcGenIns_io_npcSrc),
    .io_pc(dnpcGenIns_io_pc),
    .io_imme(dnpcGenIns_io_imme),
    .io_rd(dnpcGenIns_io_rd),
    .io_dnpc(dnpcGenIns_io_dnpc)
  );
  memData memData_ins ( // @[execute.scala 148:27]
    .io_rdata(memData_ins_io_rdata),
    .io_rdata_ext(memData_ins_io_rdata_ext),
    .io_memReadNum(memData_ins_io_memReadNum)
  );
  assign io_dataId_dIn = _T_30 ? memData_ins_io_rdata_ext : _T_29; // @[execute.scala 165:17]
  assign io_dataOut_ALUResOut = io_CSRCtrlIf_rfen ? csr_ins_io_rd : ALU_io_ALUResult; // @[execute.scala 120:24]
  assign io_dataOut_wdata = _T_14 ? io_aluRes3 : _T_13; // @[execute.scala 121:20]
  assign io_brTake = ALU_io_ALUResult[0]; // @[execute.scala 136:13]
  assign io_dnpc = _T_23[31:0]; // @[execute.scala 134:11]
  assign startTimeCnt = csr_ins_startTimeCnt_0;
  assign block1 = ALU_block1_0;
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_srcA = _T_9 ? {{32'd0}, io_pc} : _T_8; // @[execute.scala 97:15]
  assign ALU_io_srcB = _T_19 ? {{32'd0}, io_pc} : _T_18; // @[execute.scala 98:15]
  assign ALU_io_ALUCtrl = io_ALUCtrl; // @[execute.scala 99:18]
  assign ALU_block23_0 = block23;
  assign csr_ins_clock = clock;
  assign csr_ins_reset = reset;
  assign csr_ins_io_csrrwen = io_CSRCtrlIf_csrrwen; // @[execute.scala 104:22]
  assign csr_ins_io_csrswen = io_CSRCtrlIf_csrswen; // @[execute.scala 105:22]
  assign csr_ins_io_csrrsien = io_CSRCtrlIf_csrrsien; // @[execute.scala 106:23]
  assign csr_ins_io_csrrcien = io_CSRCtrlIf_csrrcien; // @[execute.scala 107:23]
  assign csr_ins_io_csrrcen = io_CSRCtrlIf_csrrcen; // @[execute.scala 108:22]
  assign csr_ins_io_csrrwien = io_CSRCtrlIf_csrrwien; // @[execute.scala 109:23]
  assign csr_ins_io_ecall = io_CSRCtrlIf_ecall; // @[execute.scala 110:20]
  assign csr_ins_io_rs1 = _T_4 ? io_aluRes3 : _T_3; // @[execute.scala 112:18]
  assign csr_ins_io_imme = io_dataId_imme[11:0]; // @[execute.scala 113:19]
  assign csr_ins_io_pc = {{32'd0}, io_pc}; // @[execute.scala 114:17]
  assign csr_ins_io_uimm = io_uimm; // @[execute.scala 115:19]
  assign csr_ins_io_mret = io_CSRCtrlIf_mepc2pc; // @[execute.scala 116:19]
  assign csr_ins_intrTimeCnt_0 = intrTimeCnt_0;
  assign csr_ins_block1_0 = block1;
  assign csr_ins_block23_0 = block23;
  assign dnpcGenIns_io_npcSrc = io_dnpcSrc; // @[execute.scala 128:24]
  assign dnpcGenIns_io_pc = io_pc; // @[execute.scala 124:20]
  assign dnpcGenIns_io_imme = io_dataId_imme[31:0]; // @[execute.scala 125:22]
  assign dnpcGenIns_io_rd = dOut1[31:0]; // @[execute.scala 127:20]
  assign memData_ins_io_rdata = io_dataOut_rdata; // @[execute.scala 150:24]
  assign memData_ins_io_memReadNum = io_memReadNum; // @[execute.scala 149:29]
endmodule
module hazard(
  input        io_regEnEXMEM,
  input  [4:0] io_rdEXMEM,
  input  [4:0] io_rs1IDEX,
  input  [4:0] io_rs2IDEX,
  input        io_regEnMEMWB,
  input  [4:0] io_rdMEMWB,
  input        io_regEnWBEND,
  input  [4:0] io_rdWBEND,
  output [1:0] io_forwardA,
  output [1:0] io_forwardB,
  input  [4:0] io_rs1IFID,
  input  [4:0] io_rs2IFID,
  input  [4:0] io_rdIDEX,
  input  [1:0] io_resSrc,
  output       io_loadHazard
);
  wire  _T = io_rdEXMEM == io_rs1IDEX; // @[hazard.scala 36:48]
  wire  _T_1 = io_regEnEXMEM & _T; // @[hazard.scala 36:35]
  wire  _T_2 = io_rs1IDEX != 5'h0; // @[hazard.scala 36:76]
  wire  forwardAOne = _T_1 & _T_2; // @[hazard.scala 36:63]
  wire  _T_3 = io_rdMEMWB == io_rs1IDEX; // @[hazard.scala 37:49]
  wire  _T_4 = io_regEnMEMWB & _T_3; // @[hazard.scala 37:35]
  wire  _T_6 = _T_4 & _T_2; // @[hazard.scala 37:64]
  wire  _T_7 = io_rdEXMEM != io_rs1IDEX; // @[hazard.scala 37:97]
  wire  _T_8 = ~io_regEnEXMEM; // @[hazard.scala 37:115]
  wire  _T_9 = _T_7 | _T_8; // @[hazard.scala 37:112]
  wire  forwardATwo = _T_6 & _T_9; // @[hazard.scala 37:84]
  wire  _T_10 = io_rdWBEND == io_rs1IDEX; // @[hazard.scala 38:51]
  wire  _T_11 = io_regEnWBEND & _T_10; // @[hazard.scala 38:37]
  wire  forwardAThree = _T_11 & _T_2; // @[hazard.scala 38:66]
  wire [1:0] _T_13 = forwardAThree ? 2'h3 : 2'h0; // @[hazard.scala 39:75]
  wire [1:0] _T_14 = forwardATwo ? 2'h1 : _T_13; // @[hazard.scala 39:47]
  wire  _T_16 = io_rdEXMEM == io_rs2IDEX; // @[hazard.scala 41:48]
  wire  _T_17 = io_regEnEXMEM & _T_16; // @[hazard.scala 41:35]
  wire  _T_18 = io_rs2IDEX != 5'h0; // @[hazard.scala 41:76]
  wire  forwardBOne = _T_17 & _T_18; // @[hazard.scala 41:63]
  wire  _T_19 = io_rdMEMWB == io_rs2IDEX; // @[hazard.scala 42:49]
  wire  _T_20 = io_regEnMEMWB & _T_19; // @[hazard.scala 42:35]
  wire  _T_22 = _T_20 & _T_18; // @[hazard.scala 42:64]
  wire  _T_23 = io_rdEXMEM != io_rs2IDEX; // @[hazard.scala 42:97]
  wire  _T_25 = _T_23 | _T_8; // @[hazard.scala 42:112]
  wire  forwardBTwo = _T_22 & _T_25; // @[hazard.scala 42:84]
  wire  _T_26 = io_rdWBEND == io_rs2IDEX; // @[hazard.scala 43:52]
  wire  _T_27 = io_regEnWBEND & _T_26; // @[hazard.scala 43:38]
  wire  forwardBThree = _T_27 & _T_18; // @[hazard.scala 43:67]
  wire [1:0] _T_29 = forwardBThree ? 2'h3 : 2'h0; // @[hazard.scala 44:75]
  wire [1:0] _T_30 = forwardBTwo ? 2'h1 : _T_29; // @[hazard.scala 44:47]
  wire  _T_32 = io_rs1IFID == io_rdIDEX; // @[hazard.scala 46:32]
  wire  _T_33 = io_rs2IFID == io_rdIDEX; // @[hazard.scala 46:59]
  wire  _T_34 = _T_32 | _T_33; // @[hazard.scala 46:46]
  wire  _T_35 = io_resSrc == 2'h2; // @[hazard.scala 46:87]
  assign io_forwardA = forwardAOne ? 2'h2 : _T_14; // @[hazard.scala 39:15]
  assign io_forwardB = forwardBOne ? 2'h2 : _T_30; // @[hazard.scala 44:15]
  assign io_loadHazard = _T_34 & _T_35; // @[hazard.scala 46:17]
endmodule
module preCell(
  input         clock,
  input         reset,
  input         io_cen,
  input         io_jump,
  input  [31:0] io_dnpcIn,
  output [31:0] io_dnpcOut,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _T = io_cen & io_jump; // @[preCell.scala 16:48]
  reg [31:0] dnpcReg; // @[Reg.scala 27:20]
  wire  takenV = dnpcReg == io_dnpcIn; // @[preCell.scala 21:24]
  reg [1:0] stateWire; // @[Reg.scala 27:20]
  wire  _T_1 = 2'h1 == stateWire; // @[Mux.scala 80:60]
  wire  _T_3 = 2'h2 == stateWire; // @[Mux.scala 80:60]
  wire  _T_5 = 2'h3 == stateWire; // @[Mux.scala 80:60]
  wire  _T_8 = stateWire == 2'h2; // @[preCell.scala 43:25]
  wire  _T_9 = stateWire == 2'h3; // @[preCell.scala 43:49]
  assign io_dnpcOut = dnpcReg; // @[preCell.scala 42:14]
  assign io_valid = _T_8 | _T_9; // @[preCell.scala 43:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dnpcReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stateWire = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      dnpcReg <= 32'h0;
    end else if (_T) begin
      dnpcReg <= io_dnpcIn;
    end
    if (reset) begin
      stateWire <= 2'h0;
    end else if (io_cen) begin
      if (_T_5) begin
        if (takenV) begin
          stateWire <= 2'h3;
        end else begin
          stateWire <= 2'h2;
        end
      end else if (_T_3) begin
        if (takenV) begin
          stateWire <= 2'h3;
        end else begin
          stateWire <= 2'h1;
        end
      end else if (_T_1) begin
        if (takenV) begin
          stateWire <= 2'h2;
        end else begin
          stateWire <= 2'h0;
        end
      end else if (takenV) begin
        stateWire <= 2'h1;
      end else begin
        stateWire <= 2'h0;
      end
    end
  end
endmodule
module preBranch(
  input         clock,
  input         reset,
  input         io_exjump,
  input  [31:0] io_ifpc,
  input  [31:0] io_expc,
  input  [31:0] io_exdpc,
  output [31:0] io_ifdnpc,
  output        io_ifjump,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  precelList_0_clock; // @[preBranch.scala 27:45]
  wire  precelList_0_reset; // @[preBranch.scala 27:45]
  wire  precelList_0_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_0_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_0_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_0_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_0_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_1_clock; // @[preBranch.scala 27:45]
  wire  precelList_1_reset; // @[preBranch.scala 27:45]
  wire  precelList_1_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_1_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_1_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_1_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_1_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_2_clock; // @[preBranch.scala 27:45]
  wire  precelList_2_reset; // @[preBranch.scala 27:45]
  wire  precelList_2_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_2_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_2_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_2_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_2_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_3_clock; // @[preBranch.scala 27:45]
  wire  precelList_3_reset; // @[preBranch.scala 27:45]
  wire  precelList_3_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_3_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_3_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_3_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_3_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_4_clock; // @[preBranch.scala 27:45]
  wire  precelList_4_reset; // @[preBranch.scala 27:45]
  wire  precelList_4_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_4_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_4_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_4_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_4_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_5_clock; // @[preBranch.scala 27:45]
  wire  precelList_5_reset; // @[preBranch.scala 27:45]
  wire  precelList_5_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_5_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_5_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_5_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_5_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_6_clock; // @[preBranch.scala 27:45]
  wire  precelList_6_reset; // @[preBranch.scala 27:45]
  wire  precelList_6_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_6_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_6_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_6_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_6_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_7_clock; // @[preBranch.scala 27:45]
  wire  precelList_7_reset; // @[preBranch.scala 27:45]
  wire  precelList_7_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_7_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_7_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_7_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_7_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_8_clock; // @[preBranch.scala 27:45]
  wire  precelList_8_reset; // @[preBranch.scala 27:45]
  wire  precelList_8_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_8_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_8_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_8_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_8_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_9_clock; // @[preBranch.scala 27:45]
  wire  precelList_9_reset; // @[preBranch.scala 27:45]
  wire  precelList_9_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_9_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_9_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_9_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_9_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_10_clock; // @[preBranch.scala 27:45]
  wire  precelList_10_reset; // @[preBranch.scala 27:45]
  wire  precelList_10_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_10_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_10_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_10_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_10_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_11_clock; // @[preBranch.scala 27:45]
  wire  precelList_11_reset; // @[preBranch.scala 27:45]
  wire  precelList_11_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_11_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_11_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_11_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_11_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_12_clock; // @[preBranch.scala 27:45]
  wire  precelList_12_reset; // @[preBranch.scala 27:45]
  wire  precelList_12_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_12_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_12_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_12_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_12_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_13_clock; // @[preBranch.scala 27:45]
  wire  precelList_13_reset; // @[preBranch.scala 27:45]
  wire  precelList_13_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_13_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_13_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_13_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_13_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_14_clock; // @[preBranch.scala 27:45]
  wire  precelList_14_reset; // @[preBranch.scala 27:45]
  wire  precelList_14_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_14_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_14_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_14_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_14_io_valid; // @[preBranch.scala 27:45]
  wire  precelList_15_clock; // @[preBranch.scala 27:45]
  wire  precelList_15_reset; // @[preBranch.scala 27:45]
  wire  precelList_15_io_cen; // @[preBranch.scala 27:45]
  wire  precelList_15_io_jump; // @[preBranch.scala 27:45]
  wire [31:0] precelList_15_io_dnpcIn; // @[preBranch.scala 27:45]
  wire [31:0] precelList_15_io_dnpcOut; // @[preBranch.scala 27:45]
  wire  precelList_15_io_valid; // @[preBranch.scala 27:45]
  wire  block = block1_0 | block23_0; // @[preBranch.scala 24:22]
  reg [31:0] pcList_0; // @[Reg.scala 27:20]
  wire  _T = io_expc == pcList_0; // @[preBranch.scala 33:27]
  reg  vList_0; // @[Reg.scala 27:20]
  wire  hitList_0 = _T & vList_0; // @[preBranch.scala 33:41]
  reg [31:0] pcList_1; // @[Reg.scala 27:20]
  wire  _T_2 = io_expc == pcList_1; // @[preBranch.scala 33:27]
  reg  vList_1; // @[Reg.scala 27:20]
  wire  hitList_1 = _T_2 & vList_1; // @[preBranch.scala 33:41]
  reg [31:0] pcList_2; // @[Reg.scala 27:20]
  wire  _T_4 = io_expc == pcList_2; // @[preBranch.scala 33:27]
  reg  vList_2; // @[Reg.scala 27:20]
  wire  hitList_2 = _T_4 & vList_2; // @[preBranch.scala 33:41]
  reg [31:0] pcList_3; // @[Reg.scala 27:20]
  wire  _T_6 = io_expc == pcList_3; // @[preBranch.scala 33:27]
  reg  vList_3; // @[Reg.scala 27:20]
  wire  hitList_3 = _T_6 & vList_3; // @[preBranch.scala 33:41]
  reg [31:0] pcList_4; // @[Reg.scala 27:20]
  wire  _T_8 = io_expc == pcList_4; // @[preBranch.scala 33:27]
  reg  vList_4; // @[Reg.scala 27:20]
  wire  hitList_4 = _T_8 & vList_4; // @[preBranch.scala 33:41]
  reg [31:0] pcList_5; // @[Reg.scala 27:20]
  wire  _T_10 = io_expc == pcList_5; // @[preBranch.scala 33:27]
  reg  vList_5; // @[Reg.scala 27:20]
  wire  hitList_5 = _T_10 & vList_5; // @[preBranch.scala 33:41]
  reg [31:0] pcList_6; // @[Reg.scala 27:20]
  wire  _T_12 = io_expc == pcList_6; // @[preBranch.scala 33:27]
  reg  vList_6; // @[Reg.scala 27:20]
  wire  hitList_6 = _T_12 & vList_6; // @[preBranch.scala 33:41]
  reg [31:0] pcList_7; // @[Reg.scala 27:20]
  wire  _T_14 = io_expc == pcList_7; // @[preBranch.scala 33:27]
  reg  vList_7; // @[Reg.scala 27:20]
  wire  hitList_7 = _T_14 & vList_7; // @[preBranch.scala 33:41]
  reg [31:0] pcList_8; // @[Reg.scala 27:20]
  wire  _T_16 = io_expc == pcList_8; // @[preBranch.scala 33:27]
  reg  vList_8; // @[Reg.scala 27:20]
  wire  hitList_8 = _T_16 & vList_8; // @[preBranch.scala 33:41]
  reg [31:0] pcList_9; // @[Reg.scala 27:20]
  wire  _T_18 = io_expc == pcList_9; // @[preBranch.scala 33:27]
  reg  vList_9; // @[Reg.scala 27:20]
  wire  hitList_9 = _T_18 & vList_9; // @[preBranch.scala 33:41]
  reg [31:0] pcList_10; // @[Reg.scala 27:20]
  wire  _T_20 = io_expc == pcList_10; // @[preBranch.scala 33:27]
  reg  vList_10; // @[Reg.scala 27:20]
  wire  hitList_10 = _T_20 & vList_10; // @[preBranch.scala 33:41]
  reg [31:0] pcList_11; // @[Reg.scala 27:20]
  wire  _T_22 = io_expc == pcList_11; // @[preBranch.scala 33:27]
  reg  vList_11; // @[Reg.scala 27:20]
  wire  hitList_11 = _T_22 & vList_11; // @[preBranch.scala 33:41]
  reg [31:0] pcList_12; // @[Reg.scala 27:20]
  wire  _T_24 = io_expc == pcList_12; // @[preBranch.scala 33:27]
  reg  vList_12; // @[Reg.scala 27:20]
  wire  hitList_12 = _T_24 & vList_12; // @[preBranch.scala 33:41]
  reg [31:0] pcList_13; // @[Reg.scala 27:20]
  wire  _T_26 = io_expc == pcList_13; // @[preBranch.scala 33:27]
  reg  vList_13; // @[Reg.scala 27:20]
  wire  hitList_13 = _T_26 & vList_13; // @[preBranch.scala 33:41]
  reg [31:0] pcList_14; // @[Reg.scala 27:20]
  wire  _T_28 = io_expc == pcList_14; // @[preBranch.scala 33:27]
  reg  vList_14; // @[Reg.scala 27:20]
  wire  hitList_14 = _T_28 & vList_14; // @[preBranch.scala 33:41]
  reg [31:0] pcList_15; // @[Reg.scala 27:20]
  wire  _T_30 = io_expc == pcList_15; // @[preBranch.scala 33:27]
  reg  vList_15; // @[Reg.scala 27:20]
  wire  hitList_15 = _T_30 & vList_15; // @[preBranch.scala 33:41]
  wire  _T_33 = hitList_0 | hitList_1; // @[preBranch.scala 35:51]
  wire  _T_34 = _T_33 | hitList_2; // @[preBranch.scala 35:51]
  wire  _T_35 = _T_34 | hitList_3; // @[preBranch.scala 35:51]
  wire  _T_36 = _T_35 | hitList_4; // @[preBranch.scala 35:51]
  wire  _T_37 = _T_36 | hitList_5; // @[preBranch.scala 35:51]
  wire  _T_38 = _T_37 | hitList_6; // @[preBranch.scala 35:51]
  wire  _T_39 = _T_38 | hitList_7; // @[preBranch.scala 35:51]
  wire  _T_40 = _T_39 | hitList_8; // @[preBranch.scala 35:51]
  wire  _T_41 = _T_40 | hitList_9; // @[preBranch.scala 35:51]
  wire  _T_42 = _T_41 | hitList_10; // @[preBranch.scala 35:51]
  wire  _T_43 = _T_42 | hitList_11; // @[preBranch.scala 35:51]
  wire  _T_44 = _T_43 | hitList_12; // @[preBranch.scala 35:51]
  wire  _T_45 = _T_44 | hitList_13; // @[preBranch.scala 35:51]
  wire  _T_46 = _T_45 | hitList_14; // @[preBranch.scala 35:51]
  wire  hit = _T_46 | hitList_15; // @[preBranch.scala 35:51]
  reg [3:0] cnt; // @[Reg.scala 27:20]
  wire [3:0] _T_48 = cnt + 4'h1; // @[preBranch.scala 38:25]
  wire  _T_49 = ~hit; // @[preBranch.scala 38:40]
  wire  _T_50 = _T_49 & io_exjump; // @[preBranch.scala 38:45]
  wire  _T_51 = ~block; // @[preBranch.scala 38:61]
  wire  _T_52 = _T_50 & _T_51; // @[preBranch.scala 38:58]
  wire  _T_54 = cnt == 4'h0; // @[preBranch.scala 44:62]
  wire  _T_55 = io_exjump & _T_54; // @[preBranch.scala 44:55]
  wire  _T_56 = hitList_0 | _T_55; // @[preBranch.scala 44:41]
  wire  _T_59 = ~hitList_0; // @[preBranch.scala 46:44]
  wire  _T_60 = _T_59 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_62 = _T_60 & _T_54; // @[preBranch.scala 46:67]
  wire  _T_64 = _T_62 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_1 = _T_64 | vList_0; // @[Reg.scala 28:19]
  wire  _T_73 = cnt == 4'h1; // @[preBranch.scala 44:62]
  wire  _T_74 = io_exjump & _T_73; // @[preBranch.scala 44:55]
  wire  _T_75 = hitList_1 | _T_74; // @[preBranch.scala 44:41]
  wire  _T_78 = ~hitList_1; // @[preBranch.scala 46:44]
  wire  _T_79 = _T_78 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_81 = _T_79 & _T_73; // @[preBranch.scala 46:67]
  wire  _T_83 = _T_81 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_3 = _T_83 | vList_1; // @[Reg.scala 28:19]
  wire  _T_92 = cnt == 4'h2; // @[preBranch.scala 44:62]
  wire  _T_93 = io_exjump & _T_92; // @[preBranch.scala 44:55]
  wire  _T_94 = hitList_2 | _T_93; // @[preBranch.scala 44:41]
  wire  _T_97 = ~hitList_2; // @[preBranch.scala 46:44]
  wire  _T_98 = _T_97 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_100 = _T_98 & _T_92; // @[preBranch.scala 46:67]
  wire  _T_102 = _T_100 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_5 = _T_102 | vList_2; // @[Reg.scala 28:19]
  wire  _T_111 = cnt == 4'h3; // @[preBranch.scala 44:62]
  wire  _T_112 = io_exjump & _T_111; // @[preBranch.scala 44:55]
  wire  _T_113 = hitList_3 | _T_112; // @[preBranch.scala 44:41]
  wire  _T_116 = ~hitList_3; // @[preBranch.scala 46:44]
  wire  _T_117 = _T_116 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_119 = _T_117 & _T_111; // @[preBranch.scala 46:67]
  wire  _T_121 = _T_119 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_7 = _T_121 | vList_3; // @[Reg.scala 28:19]
  wire  _T_130 = cnt == 4'h4; // @[preBranch.scala 44:62]
  wire  _T_131 = io_exjump & _T_130; // @[preBranch.scala 44:55]
  wire  _T_132 = hitList_4 | _T_131; // @[preBranch.scala 44:41]
  wire  _T_135 = ~hitList_4; // @[preBranch.scala 46:44]
  wire  _T_136 = _T_135 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_138 = _T_136 & _T_130; // @[preBranch.scala 46:67]
  wire  _T_140 = _T_138 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_9 = _T_140 | vList_4; // @[Reg.scala 28:19]
  wire  _T_149 = cnt == 4'h5; // @[preBranch.scala 44:62]
  wire  _T_150 = io_exjump & _T_149; // @[preBranch.scala 44:55]
  wire  _T_151 = hitList_5 | _T_150; // @[preBranch.scala 44:41]
  wire  _T_154 = ~hitList_5; // @[preBranch.scala 46:44]
  wire  _T_155 = _T_154 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_157 = _T_155 & _T_149; // @[preBranch.scala 46:67]
  wire  _T_159 = _T_157 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_11 = _T_159 | vList_5; // @[Reg.scala 28:19]
  wire  _T_168 = cnt == 4'h6; // @[preBranch.scala 44:62]
  wire  _T_169 = io_exjump & _T_168; // @[preBranch.scala 44:55]
  wire  _T_170 = hitList_6 | _T_169; // @[preBranch.scala 44:41]
  wire  _T_173 = ~hitList_6; // @[preBranch.scala 46:44]
  wire  _T_174 = _T_173 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_176 = _T_174 & _T_168; // @[preBranch.scala 46:67]
  wire  _T_178 = _T_176 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_13 = _T_178 | vList_6; // @[Reg.scala 28:19]
  wire  _T_187 = cnt == 4'h7; // @[preBranch.scala 44:62]
  wire  _T_188 = io_exjump & _T_187; // @[preBranch.scala 44:55]
  wire  _T_189 = hitList_7 | _T_188; // @[preBranch.scala 44:41]
  wire  _T_192 = ~hitList_7; // @[preBranch.scala 46:44]
  wire  _T_193 = _T_192 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_195 = _T_193 & _T_187; // @[preBranch.scala 46:67]
  wire  _T_197 = _T_195 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_15 = _T_197 | vList_7; // @[Reg.scala 28:19]
  wire  _T_206 = cnt == 4'h8; // @[preBranch.scala 44:62]
  wire  _T_207 = io_exjump & _T_206; // @[preBranch.scala 44:55]
  wire  _T_208 = hitList_8 | _T_207; // @[preBranch.scala 44:41]
  wire  _T_211 = ~hitList_8; // @[preBranch.scala 46:44]
  wire  _T_212 = _T_211 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_214 = _T_212 & _T_206; // @[preBranch.scala 46:67]
  wire  _T_216 = _T_214 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_17 = _T_216 | vList_8; // @[Reg.scala 28:19]
  wire  _T_225 = cnt == 4'h9; // @[preBranch.scala 44:62]
  wire  _T_226 = io_exjump & _T_225; // @[preBranch.scala 44:55]
  wire  _T_227 = hitList_9 | _T_226; // @[preBranch.scala 44:41]
  wire  _T_230 = ~hitList_9; // @[preBranch.scala 46:44]
  wire  _T_231 = _T_230 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_233 = _T_231 & _T_225; // @[preBranch.scala 46:67]
  wire  _T_235 = _T_233 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_19 = _T_235 | vList_9; // @[Reg.scala 28:19]
  wire  _T_244 = cnt == 4'ha; // @[preBranch.scala 44:62]
  wire  _T_245 = io_exjump & _T_244; // @[preBranch.scala 44:55]
  wire  _T_246 = hitList_10 | _T_245; // @[preBranch.scala 44:41]
  wire  _T_249 = ~hitList_10; // @[preBranch.scala 46:44]
  wire  _T_250 = _T_249 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_252 = _T_250 & _T_244; // @[preBranch.scala 46:67]
  wire  _T_254 = _T_252 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_21 = _T_254 | vList_10; // @[Reg.scala 28:19]
  wire  _T_263 = cnt == 4'hb; // @[preBranch.scala 44:62]
  wire  _T_264 = io_exjump & _T_263; // @[preBranch.scala 44:55]
  wire  _T_265 = hitList_11 | _T_264; // @[preBranch.scala 44:41]
  wire  _T_268 = ~hitList_11; // @[preBranch.scala 46:44]
  wire  _T_269 = _T_268 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_271 = _T_269 & _T_263; // @[preBranch.scala 46:67]
  wire  _T_273 = _T_271 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_23 = _T_273 | vList_11; // @[Reg.scala 28:19]
  wire  _T_282 = cnt == 4'hc; // @[preBranch.scala 44:62]
  wire  _T_283 = io_exjump & _T_282; // @[preBranch.scala 44:55]
  wire  _T_284 = hitList_12 | _T_283; // @[preBranch.scala 44:41]
  wire  _T_287 = ~hitList_12; // @[preBranch.scala 46:44]
  wire  _T_288 = _T_287 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_290 = _T_288 & _T_282; // @[preBranch.scala 46:67]
  wire  _T_292 = _T_290 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_25 = _T_292 | vList_12; // @[Reg.scala 28:19]
  wire  _T_301 = cnt == 4'hd; // @[preBranch.scala 44:62]
  wire  _T_302 = io_exjump & _T_301; // @[preBranch.scala 44:55]
  wire  _T_303 = hitList_13 | _T_302; // @[preBranch.scala 44:41]
  wire  _T_306 = ~hitList_13; // @[preBranch.scala 46:44]
  wire  _T_307 = _T_306 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_309 = _T_307 & _T_301; // @[preBranch.scala 46:67]
  wire  _T_311 = _T_309 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_27 = _T_311 | vList_13; // @[Reg.scala 28:19]
  wire  _T_320 = cnt == 4'he; // @[preBranch.scala 44:62]
  wire  _T_321 = io_exjump & _T_320; // @[preBranch.scala 44:55]
  wire  _T_322 = hitList_14 | _T_321; // @[preBranch.scala 44:41]
  wire  _T_325 = ~hitList_14; // @[preBranch.scala 46:44]
  wire  _T_326 = _T_325 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_328 = _T_326 & _T_320; // @[preBranch.scala 46:67]
  wire  _T_330 = _T_328 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_29 = _T_330 | vList_14; // @[Reg.scala 28:19]
  wire  _T_339 = cnt == 4'hf; // @[preBranch.scala 44:62]
  wire  _T_340 = io_exjump & _T_339; // @[preBranch.scala 44:55]
  wire  _T_341 = hitList_15 | _T_340; // @[preBranch.scala 44:41]
  wire  _T_344 = ~hitList_15; // @[preBranch.scala 46:44]
  wire  _T_345 = _T_344 & io_exjump; // @[preBranch.scala 46:55]
  wire  _T_347 = _T_345 & _T_339; // @[preBranch.scala 46:67]
  wire  _T_349 = _T_347 & _T_51; // @[preBranch.scala 46:82]
  wire  _GEN_31 = _T_349 | vList_15; // @[Reg.scala 28:19]
  wire  _T_358 = io_ifpc == pcList_0; // @[preBranch.scala 55:29]
  wire  hitIfList_0 = _T_358 & vList_0; // @[preBranch.scala 55:43]
  wire  _T_360 = io_ifpc == pcList_1; // @[preBranch.scala 55:29]
  wire  hitIfList_1 = _T_360 & vList_1; // @[preBranch.scala 55:43]
  wire  _T_362 = io_ifpc == pcList_2; // @[preBranch.scala 55:29]
  wire  hitIfList_2 = _T_362 & vList_2; // @[preBranch.scala 55:43]
  wire  _T_364 = io_ifpc == pcList_3; // @[preBranch.scala 55:29]
  wire  hitIfList_3 = _T_364 & vList_3; // @[preBranch.scala 55:43]
  wire  _T_366 = io_ifpc == pcList_4; // @[preBranch.scala 55:29]
  wire  hitIfList_4 = _T_366 & vList_4; // @[preBranch.scala 55:43]
  wire  _T_368 = io_ifpc == pcList_5; // @[preBranch.scala 55:29]
  wire  hitIfList_5 = _T_368 & vList_5; // @[preBranch.scala 55:43]
  wire  _T_370 = io_ifpc == pcList_6; // @[preBranch.scala 55:29]
  wire  hitIfList_6 = _T_370 & vList_6; // @[preBranch.scala 55:43]
  wire  _T_372 = io_ifpc == pcList_7; // @[preBranch.scala 55:29]
  wire  hitIfList_7 = _T_372 & vList_7; // @[preBranch.scala 55:43]
  wire  _T_374 = io_ifpc == pcList_8; // @[preBranch.scala 55:29]
  wire  hitIfList_8 = _T_374 & vList_8; // @[preBranch.scala 55:43]
  wire  _T_376 = io_ifpc == pcList_9; // @[preBranch.scala 55:29]
  wire  hitIfList_9 = _T_376 & vList_9; // @[preBranch.scala 55:43]
  wire  _T_378 = io_ifpc == pcList_10; // @[preBranch.scala 55:29]
  wire  hitIfList_10 = _T_378 & vList_10; // @[preBranch.scala 55:43]
  wire  _T_380 = io_ifpc == pcList_11; // @[preBranch.scala 55:29]
  wire  hitIfList_11 = _T_380 & vList_11; // @[preBranch.scala 55:43]
  wire  _T_382 = io_ifpc == pcList_12; // @[preBranch.scala 55:29]
  wire  hitIfList_12 = _T_382 & vList_12; // @[preBranch.scala 55:43]
  wire  _T_384 = io_ifpc == pcList_13; // @[preBranch.scala 55:29]
  wire  hitIfList_13 = _T_384 & vList_13; // @[preBranch.scala 55:43]
  wire  _T_386 = io_ifpc == pcList_14; // @[preBranch.scala 55:29]
  wire  hitIfList_14 = _T_386 & vList_14; // @[preBranch.scala 55:43]
  wire  _T_388 = io_ifpc == pcList_15; // @[preBranch.scala 55:29]
  wire  hitIfList_15 = _T_388 & vList_15; // @[preBranch.scala 55:43]
  wire  _T_391 = hitIfList_0 | hitIfList_1; // @[preBranch.scala 58:55]
  wire  _T_392 = _T_391 | hitIfList_2; // @[preBranch.scala 58:55]
  wire  _T_393 = _T_392 | hitIfList_3; // @[preBranch.scala 58:55]
  wire  _T_394 = _T_393 | hitIfList_4; // @[preBranch.scala 58:55]
  wire  _T_395 = _T_394 | hitIfList_5; // @[preBranch.scala 58:55]
  wire  _T_396 = _T_395 | hitIfList_6; // @[preBranch.scala 58:55]
  wire  _T_397 = _T_396 | hitIfList_7; // @[preBranch.scala 58:55]
  wire  _T_398 = _T_397 | hitIfList_8; // @[preBranch.scala 58:55]
  wire  _T_399 = _T_398 | hitIfList_9; // @[preBranch.scala 58:55]
  wire  _T_400 = _T_399 | hitIfList_10; // @[preBranch.scala 58:55]
  wire  _T_401 = _T_400 | hitIfList_11; // @[preBranch.scala 58:55]
  wire  _T_402 = _T_401 | hitIfList_12; // @[preBranch.scala 58:55]
  wire  _T_403 = _T_402 | hitIfList_13; // @[preBranch.scala 58:55]
  wire  _T_404 = _T_403 | hitIfList_14; // @[preBranch.scala 58:55]
  wire  hitif = _T_404 | hitIfList_15; // @[preBranch.scala 58:55]
  wire  _T_405 = ~hitif; // @[preBranch.scala 64:5]
  wire  _T_406 = hitIfList_0 & precelList_0_io_valid; // @[Mux.scala 27:72]
  wire  _T_407 = hitIfList_1 & precelList_1_io_valid; // @[Mux.scala 27:72]
  wire  _T_408 = hitIfList_2 & precelList_2_io_valid; // @[Mux.scala 27:72]
  wire  _T_409 = hitIfList_3 & precelList_3_io_valid; // @[Mux.scala 27:72]
  wire  _T_410 = hitIfList_4 & precelList_4_io_valid; // @[Mux.scala 27:72]
  wire  _T_411 = hitIfList_5 & precelList_5_io_valid; // @[Mux.scala 27:72]
  wire  _T_412 = hitIfList_6 & precelList_6_io_valid; // @[Mux.scala 27:72]
  wire  _T_413 = hitIfList_7 & precelList_7_io_valid; // @[Mux.scala 27:72]
  wire  _T_414 = hitIfList_8 & precelList_8_io_valid; // @[Mux.scala 27:72]
  wire  _T_415 = hitIfList_9 & precelList_9_io_valid; // @[Mux.scala 27:72]
  wire  _T_416 = hitIfList_10 & precelList_10_io_valid; // @[Mux.scala 27:72]
  wire  _T_417 = hitIfList_11 & precelList_11_io_valid; // @[Mux.scala 27:72]
  wire  _T_418 = hitIfList_12 & precelList_12_io_valid; // @[Mux.scala 27:72]
  wire  _T_419 = hitIfList_13 & precelList_13_io_valid; // @[Mux.scala 27:72]
  wire  _T_420 = hitIfList_14 & precelList_14_io_valid; // @[Mux.scala 27:72]
  wire  _T_421 = hitIfList_15 & precelList_15_io_valid; // @[Mux.scala 27:72]
  wire  _T_422 = _T_406 | _T_407; // @[Mux.scala 27:72]
  wire  _T_423 = _T_422 | _T_408; // @[Mux.scala 27:72]
  wire  _T_424 = _T_423 | _T_409; // @[Mux.scala 27:72]
  wire  _T_425 = _T_424 | _T_410; // @[Mux.scala 27:72]
  wire  _T_426 = _T_425 | _T_411; // @[Mux.scala 27:72]
  wire  _T_427 = _T_426 | _T_412; // @[Mux.scala 27:72]
  wire  _T_428 = _T_427 | _T_413; // @[Mux.scala 27:72]
  wire  _T_429 = _T_428 | _T_414; // @[Mux.scala 27:72]
  wire  _T_430 = _T_429 | _T_415; // @[Mux.scala 27:72]
  wire  _T_431 = _T_430 | _T_416; // @[Mux.scala 27:72]
  wire  _T_432 = _T_431 | _T_417; // @[Mux.scala 27:72]
  wire  _T_433 = _T_432 | _T_418; // @[Mux.scala 27:72]
  wire  _T_434 = _T_433 | _T_419; // @[Mux.scala 27:72]
  wire  _T_435 = _T_434 | _T_420; // @[Mux.scala 27:72]
  wire  _T_436 = _T_435 | _T_421; // @[Mux.scala 27:72]
  wire [31:0] _T_440 = hitIfList_0 ? precelList_0_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_441 = hitIfList_1 ? precelList_1_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_442 = hitIfList_2 ? precelList_2_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_443 = hitIfList_3 ? precelList_3_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_444 = hitIfList_4 ? precelList_4_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_445 = hitIfList_5 ? precelList_5_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_446 = hitIfList_6 ? precelList_6_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_447 = hitIfList_7 ? precelList_7_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_448 = hitIfList_8 ? precelList_8_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_449 = hitIfList_9 ? precelList_9_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_450 = hitIfList_10 ? precelList_10_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_451 = hitIfList_11 ? precelList_11_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_452 = hitIfList_12 ? precelList_12_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_453 = hitIfList_13 ? precelList_13_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_454 = hitIfList_14 ? precelList_14_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_455 = hitIfList_15 ? precelList_15_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_456 = _T_440 | _T_441; // @[Mux.scala 27:72]
  wire [31:0] _T_457 = _T_456 | _T_442; // @[Mux.scala 27:72]
  wire [31:0] _T_458 = _T_457 | _T_443; // @[Mux.scala 27:72]
  wire [31:0] _T_459 = _T_458 | _T_444; // @[Mux.scala 27:72]
  wire [31:0] _T_460 = _T_459 | _T_445; // @[Mux.scala 27:72]
  wire [31:0] _T_461 = _T_460 | _T_446; // @[Mux.scala 27:72]
  wire [31:0] _T_462 = _T_461 | _T_447; // @[Mux.scala 27:72]
  wire [31:0] _T_463 = _T_462 | _T_448; // @[Mux.scala 27:72]
  wire [31:0] _T_464 = _T_463 | _T_449; // @[Mux.scala 27:72]
  wire [31:0] _T_465 = _T_464 | _T_450; // @[Mux.scala 27:72]
  wire [31:0] _T_466 = _T_465 | _T_451; // @[Mux.scala 27:72]
  wire [31:0] _T_467 = _T_466 | _T_452; // @[Mux.scala 27:72]
  wire [31:0] _T_468 = _T_467 | _T_453; // @[Mux.scala 27:72]
  wire [31:0] _T_469 = _T_468 | _T_454; // @[Mux.scala 27:72]
  wire [31:0] _T_470 = _T_469 | _T_455; // @[Mux.scala 27:72]
  preCell precelList_0 ( // @[preBranch.scala 27:45]
    .clock(precelList_0_clock),
    .reset(precelList_0_reset),
    .io_cen(precelList_0_io_cen),
    .io_jump(precelList_0_io_jump),
    .io_dnpcIn(precelList_0_io_dnpcIn),
    .io_dnpcOut(precelList_0_io_dnpcOut),
    .io_valid(precelList_0_io_valid)
  );
  preCell precelList_1 ( // @[preBranch.scala 27:45]
    .clock(precelList_1_clock),
    .reset(precelList_1_reset),
    .io_cen(precelList_1_io_cen),
    .io_jump(precelList_1_io_jump),
    .io_dnpcIn(precelList_1_io_dnpcIn),
    .io_dnpcOut(precelList_1_io_dnpcOut),
    .io_valid(precelList_1_io_valid)
  );
  preCell precelList_2 ( // @[preBranch.scala 27:45]
    .clock(precelList_2_clock),
    .reset(precelList_2_reset),
    .io_cen(precelList_2_io_cen),
    .io_jump(precelList_2_io_jump),
    .io_dnpcIn(precelList_2_io_dnpcIn),
    .io_dnpcOut(precelList_2_io_dnpcOut),
    .io_valid(precelList_2_io_valid)
  );
  preCell precelList_3 ( // @[preBranch.scala 27:45]
    .clock(precelList_3_clock),
    .reset(precelList_3_reset),
    .io_cen(precelList_3_io_cen),
    .io_jump(precelList_3_io_jump),
    .io_dnpcIn(precelList_3_io_dnpcIn),
    .io_dnpcOut(precelList_3_io_dnpcOut),
    .io_valid(precelList_3_io_valid)
  );
  preCell precelList_4 ( // @[preBranch.scala 27:45]
    .clock(precelList_4_clock),
    .reset(precelList_4_reset),
    .io_cen(precelList_4_io_cen),
    .io_jump(precelList_4_io_jump),
    .io_dnpcIn(precelList_4_io_dnpcIn),
    .io_dnpcOut(precelList_4_io_dnpcOut),
    .io_valid(precelList_4_io_valid)
  );
  preCell precelList_5 ( // @[preBranch.scala 27:45]
    .clock(precelList_5_clock),
    .reset(precelList_5_reset),
    .io_cen(precelList_5_io_cen),
    .io_jump(precelList_5_io_jump),
    .io_dnpcIn(precelList_5_io_dnpcIn),
    .io_dnpcOut(precelList_5_io_dnpcOut),
    .io_valid(precelList_5_io_valid)
  );
  preCell precelList_6 ( // @[preBranch.scala 27:45]
    .clock(precelList_6_clock),
    .reset(precelList_6_reset),
    .io_cen(precelList_6_io_cen),
    .io_jump(precelList_6_io_jump),
    .io_dnpcIn(precelList_6_io_dnpcIn),
    .io_dnpcOut(precelList_6_io_dnpcOut),
    .io_valid(precelList_6_io_valid)
  );
  preCell precelList_7 ( // @[preBranch.scala 27:45]
    .clock(precelList_7_clock),
    .reset(precelList_7_reset),
    .io_cen(precelList_7_io_cen),
    .io_jump(precelList_7_io_jump),
    .io_dnpcIn(precelList_7_io_dnpcIn),
    .io_dnpcOut(precelList_7_io_dnpcOut),
    .io_valid(precelList_7_io_valid)
  );
  preCell precelList_8 ( // @[preBranch.scala 27:45]
    .clock(precelList_8_clock),
    .reset(precelList_8_reset),
    .io_cen(precelList_8_io_cen),
    .io_jump(precelList_8_io_jump),
    .io_dnpcIn(precelList_8_io_dnpcIn),
    .io_dnpcOut(precelList_8_io_dnpcOut),
    .io_valid(precelList_8_io_valid)
  );
  preCell precelList_9 ( // @[preBranch.scala 27:45]
    .clock(precelList_9_clock),
    .reset(precelList_9_reset),
    .io_cen(precelList_9_io_cen),
    .io_jump(precelList_9_io_jump),
    .io_dnpcIn(precelList_9_io_dnpcIn),
    .io_dnpcOut(precelList_9_io_dnpcOut),
    .io_valid(precelList_9_io_valid)
  );
  preCell precelList_10 ( // @[preBranch.scala 27:45]
    .clock(precelList_10_clock),
    .reset(precelList_10_reset),
    .io_cen(precelList_10_io_cen),
    .io_jump(precelList_10_io_jump),
    .io_dnpcIn(precelList_10_io_dnpcIn),
    .io_dnpcOut(precelList_10_io_dnpcOut),
    .io_valid(precelList_10_io_valid)
  );
  preCell precelList_11 ( // @[preBranch.scala 27:45]
    .clock(precelList_11_clock),
    .reset(precelList_11_reset),
    .io_cen(precelList_11_io_cen),
    .io_jump(precelList_11_io_jump),
    .io_dnpcIn(precelList_11_io_dnpcIn),
    .io_dnpcOut(precelList_11_io_dnpcOut),
    .io_valid(precelList_11_io_valid)
  );
  preCell precelList_12 ( // @[preBranch.scala 27:45]
    .clock(precelList_12_clock),
    .reset(precelList_12_reset),
    .io_cen(precelList_12_io_cen),
    .io_jump(precelList_12_io_jump),
    .io_dnpcIn(precelList_12_io_dnpcIn),
    .io_dnpcOut(precelList_12_io_dnpcOut),
    .io_valid(precelList_12_io_valid)
  );
  preCell precelList_13 ( // @[preBranch.scala 27:45]
    .clock(precelList_13_clock),
    .reset(precelList_13_reset),
    .io_cen(precelList_13_io_cen),
    .io_jump(precelList_13_io_jump),
    .io_dnpcIn(precelList_13_io_dnpcIn),
    .io_dnpcOut(precelList_13_io_dnpcOut),
    .io_valid(precelList_13_io_valid)
  );
  preCell precelList_14 ( // @[preBranch.scala 27:45]
    .clock(precelList_14_clock),
    .reset(precelList_14_reset),
    .io_cen(precelList_14_io_cen),
    .io_jump(precelList_14_io_jump),
    .io_dnpcIn(precelList_14_io_dnpcIn),
    .io_dnpcOut(precelList_14_io_dnpcOut),
    .io_valid(precelList_14_io_valid)
  );
  preCell precelList_15 ( // @[preBranch.scala 27:45]
    .clock(precelList_15_clock),
    .reset(precelList_15_reset),
    .io_cen(precelList_15_io_cen),
    .io_jump(precelList_15_io_jump),
    .io_dnpcIn(precelList_15_io_dnpcIn),
    .io_dnpcOut(precelList_15_io_dnpcOut),
    .io_valid(precelList_15_io_valid)
  );
  assign io_ifdnpc = _T_405 ? 32'h0 : _T_470; // @[preBranch.scala 75:13]
  assign io_ifjump = _T_405 ? 1'h0 : _T_436; // @[preBranch.scala 63:13]
  assign precelList_0_clock = clock;
  assign precelList_0_reset = reset;
  assign precelList_0_io_cen = _T_56 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_0_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_0_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_1_clock = clock;
  assign precelList_1_reset = reset;
  assign precelList_1_io_cen = _T_75 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_1_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_1_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_2_clock = clock;
  assign precelList_2_reset = reset;
  assign precelList_2_io_cen = _T_94 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_2_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_2_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_3_clock = clock;
  assign precelList_3_reset = reset;
  assign precelList_3_io_cen = _T_113 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_3_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_3_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_4_clock = clock;
  assign precelList_4_reset = reset;
  assign precelList_4_io_cen = _T_132 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_4_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_4_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_5_clock = clock;
  assign precelList_5_reset = reset;
  assign precelList_5_io_cen = _T_151 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_5_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_5_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_6_clock = clock;
  assign precelList_6_reset = reset;
  assign precelList_6_io_cen = _T_170 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_6_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_6_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_7_clock = clock;
  assign precelList_7_reset = reset;
  assign precelList_7_io_cen = _T_189 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_7_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_7_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_8_clock = clock;
  assign precelList_8_reset = reset;
  assign precelList_8_io_cen = _T_208 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_8_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_8_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_9_clock = clock;
  assign precelList_9_reset = reset;
  assign precelList_9_io_cen = _T_227 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_9_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_9_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_10_clock = clock;
  assign precelList_10_reset = reset;
  assign precelList_10_io_cen = _T_246 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_10_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_10_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_11_clock = clock;
  assign precelList_11_reset = reset;
  assign precelList_11_io_cen = _T_265 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_11_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_11_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_12_clock = clock;
  assign precelList_12_reset = reset;
  assign precelList_12_io_cen = _T_284 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_12_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_12_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_13_clock = clock;
  assign precelList_13_reset = reset;
  assign precelList_13_io_cen = _T_303 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_13_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_13_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_14_clock = clock;
  assign precelList_14_reset = reset;
  assign precelList_14_io_cen = _T_322 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_14_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_14_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
  assign precelList_15_clock = clock;
  assign precelList_15_reset = reset;
  assign precelList_15_io_cen = _T_341 & _T_51; // @[preBranch.scala 44:26]
  assign precelList_15_io_jump = io_exjump; // @[preBranch.scala 42:27]
  assign precelList_15_io_dnpcIn = io_exdpc; // @[preBranch.scala 43:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcList_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  vList_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pcList_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  vList_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pcList_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vList_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pcList_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  vList_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pcList_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  vList_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pcList_5 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  vList_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pcList_6 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  vList_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pcList_7 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  vList_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pcList_8 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  vList_8 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pcList_9 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  vList_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pcList_10 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  vList_10 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pcList_11 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  vList_11 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  pcList_12 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  vList_12 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pcList_13 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  vList_13 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pcList_14 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  vList_14 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pcList_15 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  vList_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cnt = _RAND_32[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pcList_0 <= 32'h0;
    end else if (_T_64) begin
      pcList_0 <= io_expc;
    end
    if (reset) begin
      vList_0 <= 1'h0;
    end else begin
      vList_0 <= _GEN_1;
    end
    if (reset) begin
      pcList_1 <= 32'h0;
    end else if (_T_83) begin
      pcList_1 <= io_expc;
    end
    if (reset) begin
      vList_1 <= 1'h0;
    end else begin
      vList_1 <= _GEN_3;
    end
    if (reset) begin
      pcList_2 <= 32'h0;
    end else if (_T_102) begin
      pcList_2 <= io_expc;
    end
    if (reset) begin
      vList_2 <= 1'h0;
    end else begin
      vList_2 <= _GEN_5;
    end
    if (reset) begin
      pcList_3 <= 32'h0;
    end else if (_T_121) begin
      pcList_3 <= io_expc;
    end
    if (reset) begin
      vList_3 <= 1'h0;
    end else begin
      vList_3 <= _GEN_7;
    end
    if (reset) begin
      pcList_4 <= 32'h0;
    end else if (_T_140) begin
      pcList_4 <= io_expc;
    end
    if (reset) begin
      vList_4 <= 1'h0;
    end else begin
      vList_4 <= _GEN_9;
    end
    if (reset) begin
      pcList_5 <= 32'h0;
    end else if (_T_159) begin
      pcList_5 <= io_expc;
    end
    if (reset) begin
      vList_5 <= 1'h0;
    end else begin
      vList_5 <= _GEN_11;
    end
    if (reset) begin
      pcList_6 <= 32'h0;
    end else if (_T_178) begin
      pcList_6 <= io_expc;
    end
    if (reset) begin
      vList_6 <= 1'h0;
    end else begin
      vList_6 <= _GEN_13;
    end
    if (reset) begin
      pcList_7 <= 32'h0;
    end else if (_T_197) begin
      pcList_7 <= io_expc;
    end
    if (reset) begin
      vList_7 <= 1'h0;
    end else begin
      vList_7 <= _GEN_15;
    end
    if (reset) begin
      pcList_8 <= 32'h0;
    end else if (_T_216) begin
      pcList_8 <= io_expc;
    end
    if (reset) begin
      vList_8 <= 1'h0;
    end else begin
      vList_8 <= _GEN_17;
    end
    if (reset) begin
      pcList_9 <= 32'h0;
    end else if (_T_235) begin
      pcList_9 <= io_expc;
    end
    if (reset) begin
      vList_9 <= 1'h0;
    end else begin
      vList_9 <= _GEN_19;
    end
    if (reset) begin
      pcList_10 <= 32'h0;
    end else if (_T_254) begin
      pcList_10 <= io_expc;
    end
    if (reset) begin
      vList_10 <= 1'h0;
    end else begin
      vList_10 <= _GEN_21;
    end
    if (reset) begin
      pcList_11 <= 32'h0;
    end else if (_T_273) begin
      pcList_11 <= io_expc;
    end
    if (reset) begin
      vList_11 <= 1'h0;
    end else begin
      vList_11 <= _GEN_23;
    end
    if (reset) begin
      pcList_12 <= 32'h0;
    end else if (_T_292) begin
      pcList_12 <= io_expc;
    end
    if (reset) begin
      vList_12 <= 1'h0;
    end else begin
      vList_12 <= _GEN_25;
    end
    if (reset) begin
      pcList_13 <= 32'h0;
    end else if (_T_311) begin
      pcList_13 <= io_expc;
    end
    if (reset) begin
      vList_13 <= 1'h0;
    end else begin
      vList_13 <= _GEN_27;
    end
    if (reset) begin
      pcList_14 <= 32'h0;
    end else if (_T_330) begin
      pcList_14 <= io_expc;
    end
    if (reset) begin
      vList_14 <= 1'h0;
    end else begin
      vList_14 <= _GEN_29;
    end
    if (reset) begin
      pcList_15 <= 32'h0;
    end else if (_T_349) begin
      pcList_15 <= io_expc;
    end
    if (reset) begin
      vList_15 <= 1'h0;
    end else begin
      vList_15 <= _GEN_31;
    end
    if (reset) begin
      cnt <= 4'h0;
    end else if (_T_52) begin
      cnt <= _T_48;
    end
  end
endmodule
module memVGen(
  input  [31:0] io_inst,
  output        io_valid
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memVGen.scala 20:45]
  wire  _T_1 = 32'h23 == _T; // @[memVGen.scala 20:45]
  wire  _T_3 = 32'h2023 == _T; // @[memVGen.scala 20:45]
  wire  _T_5 = 32'h3023 == _T; // @[memVGen.scala 20:45]
  wire  _T_7 = 32'h1023 == _T; // @[memVGen.scala 20:45]
  wire  _T_9 = 32'h3003 == _T; // @[memVGen.scala 26:27]
  wire  _T_11 = 32'h4003 == _T; // @[memVGen.scala 27:27]
  wire  _T_13 = 32'h1003 == _T; // @[memVGen.scala 28:27]
  wire  _T_15 = 32'h2003 == _T; // @[memVGen.scala 29:27]
  wire  _T_19 = 32'h5003 == _T; // @[memVGen.scala 31:27]
  wire  _T_21 = 32'h3 == _T; // @[memVGen.scala 32:27]
  wire  _T_23 = 32'h6003 == _T; // @[memVGen.scala 33:27]
  wire  _T_25 = _T_21 | _T_23; // @[Mux.scala 98:16]
  wire  _T_26 = _T_19 | _T_25; // @[Mux.scala 98:16]
  wire  _T_27 = _T_9 | _T_26; // @[Mux.scala 98:16]
  wire  _T_28 = _T_15 | _T_27; // @[Mux.scala 98:16]
  wire  _T_29 = _T_13 | _T_28; // @[Mux.scala 98:16]
  wire  _T_30 = _T_11 | _T_29; // @[Mux.scala 98:16]
  wire  _T_31 = _T_9 | _T_30; // @[Mux.scala 98:16]
  wire  _T_32 = _T_7 | _T_31; // @[Mux.scala 98:16]
  wire  _T_33 = _T_5 | _T_32; // @[Mux.scala 98:16]
  wire  _T_34 = _T_3 | _T_33; // @[Mux.scala 98:16]
  assign io_valid = _T_1 | _T_34; // @[memVGen.scala 36:12]
endmodule
module ALUCtrl(
  input  [31:0] io_inst,
  output [4:0]  io_ALUCtrl
);
  wire [31:0] _T = io_inst & 32'h707f; // @[ALUCtrl.scala 74:49]
  wire  _T_1 = 32'h23 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_3 = 32'h2023 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_5 = 32'h3023 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_7 = 32'h1023 == _T; // @[ALUCtrl.scala 74:49]
  wire [31:0] _T_8 = io_inst & 32'h7f; // @[ALUCtrl.scala 79:31]
  wire  _T_9 = 32'h17 == _T_8; // @[ALUCtrl.scala 79:31]
  wire  _T_11 = 32'h37 == _T_8; // @[ALUCtrl.scala 80:31]
  wire  _T_13 = 32'h13 == _T; // @[ALUCtrl.scala 81:31]
  wire  _T_15 = 32'h67 == _T; // @[ALUCtrl.scala 82:31]
  wire  _T_17 = 32'h3003 == _T; // @[ALUCtrl.scala 83:31]
  wire  _T_19 = 32'h4003 == _T; // @[ALUCtrl.scala 84:31]
  wire  _T_21 = 32'h3013 == _T; // @[ALUCtrl.scala 85:31]
  wire [31:0] _T_22 = io_inst & 32'hfe00707f; // @[ALUCtrl.scala 86:31]
  wire  _T_23 = 32'h501b == _T_22; // @[ALUCtrl.scala 86:31]
  wire [31:0] _T_24 = io_inst & 32'hfc00707f; // @[ALUCtrl.scala 87:31]
  wire  _T_25 = 32'h1013 == _T_24; // @[ALUCtrl.scala 87:31]
  wire  _T_27 = 32'h7013 == _T; // @[ALUCtrl.scala 88:31]
  wire  _T_29 = 32'h4013 == _T; // @[ALUCtrl.scala 89:31]
  wire  _T_31 = 32'h1b == _T; // @[ALUCtrl.scala 90:31]
  wire  _T_33 = 32'h5013 == _T_24; // @[ALUCtrl.scala 91:31]
  wire  _T_35 = 32'h101b == _T_22; // @[ALUCtrl.scala 92:31]
  wire  _T_37 = 32'h4000501b == _T_22; // @[ALUCtrl.scala 93:31]
  wire  _T_39 = 32'h40005013 == _T_24; // @[ALUCtrl.scala 94:31]
  wire  _T_41 = 32'h1003 == _T; // @[ALUCtrl.scala 95:31]
  wire  _T_43 = 32'h2003 == _T; // @[ALUCtrl.scala 96:31]
  wire  _T_47 = 32'h5003 == _T; // @[ALUCtrl.scala 98:31]
  wire  _T_49 = 32'h6003 == _T; // @[ALUCtrl.scala 99:31]
  wire  _T_51 = 32'h3 == _T; // @[ALUCtrl.scala 100:31]
  wire  _T_53 = 32'h6013 == _T; // @[ALUCtrl.scala 101:31]
  wire  _T_55 = 32'h3033 == _T_22; // @[ALUCtrl.scala 102:31]
  wire  _T_57 = 32'h3b == _T_22; // @[ALUCtrl.scala 103:31]
  wire  _T_59 = 32'h4000003b == _T_22; // @[ALUCtrl.scala 104:31]
  wire  _T_61 = 32'h7033 == _T_22; // @[ALUCtrl.scala 105:31]
  wire  _T_63 = 32'h33 == _T_22; // @[ALUCtrl.scala 106:31]
  wire  _T_65 = 32'h200503b == _T_22; // @[ALUCtrl.scala 107:31]
  wire  _T_67 = 32'h200703b == _T_22; // @[ALUCtrl.scala 108:31]
  wire  _T_69 = 32'h40000033 == _T_22; // @[ALUCtrl.scala 109:31]
  wire  _T_71 = 32'h200003b == _T_22; // @[ALUCtrl.scala 110:31]
  wire  _T_73 = 32'h200603b == _T_22; // @[ALUCtrl.scala 111:31]
  wire  _T_75 = 32'h200403b == _T_22; // @[ALUCtrl.scala 112:31]
  wire  _T_77 = 32'h2000033 == _T_22; // @[ALUCtrl.scala 113:31]
  wire  _T_79 = 32'h6033 == _T_22; // @[ALUCtrl.scala 114:31]
  wire  _T_81 = 32'h103b == _T_22; // @[ALUCtrl.scala 115:31]
  wire  _T_83 = 32'h4000503b == _T_22; // @[ALUCtrl.scala 116:31]
  wire  _T_85 = 32'h503b == _T_22; // @[ALUCtrl.scala 117:31]
  wire  _T_87 = 32'h2033 == _T_22; // @[ALUCtrl.scala 118:31]
  wire  _T_89 = 32'h2005033 == _T_22; // @[ALUCtrl.scala 119:31]
  wire  _T_91 = 32'h4033 == _T_22; // @[ALUCtrl.scala 120:31]
  wire  _T_93 = 32'h2006033 == _T_22; // @[ALUCtrl.scala 121:31]
  wire  _T_95 = 32'h2004033 == _T_22; // @[ALUCtrl.scala 122:31]
  wire  _T_97 = 32'h1033 == _T_22; // @[ALUCtrl.scala 123:31]
  wire  _T_99 = 32'h63 == _T; // @[ALUCtrl.scala 124:31]
  wire  _T_101 = 32'h6063 == _T; // @[ALUCtrl.scala 125:31]
  wire  _T_103 = 32'h7063 == _T; // @[ALUCtrl.scala 126:31]
  wire  _T_105 = 32'h4063 == _T; // @[ALUCtrl.scala 127:31]
  wire  _T_107 = 32'h5063 == _T; // @[ALUCtrl.scala 128:31]
  wire  _T_109 = 32'h1063 == _T; // @[ALUCtrl.scala 129:31]
  wire  _T_111 = 32'h2007033 == _T_22; // @[ALUCtrl.scala 130:31]
  wire  _T_113 = 32'h5033 == _T_22; // @[ALUCtrl.scala 131:31]
  wire [4:0] _T_114 = _T_113 ? 5'h8 : 5'h1f; // @[Mux.scala 98:16]
  wire [4:0] _T_115 = _T_111 ? 5'h1d : _T_114; // @[Mux.scala 98:16]
  wire [4:0] _T_116 = _T_109 ? 5'hb : _T_115; // @[Mux.scala 98:16]
  wire [4:0] _T_117 = _T_107 ? 5'h1c : _T_116; // @[Mux.scala 98:16]
  wire [4:0] _T_118 = _T_105 ? 5'h5 : _T_117; // @[Mux.scala 98:16]
  wire [4:0] _T_119 = _T_103 ? 5'h1b : _T_118; // @[Mux.scala 98:16]
  wire [4:0] _T_120 = _T_101 ? 5'h7 : _T_119; // @[Mux.scala 98:16]
  wire [4:0] _T_121 = _T_99 ? 5'h1a : _T_120; // @[Mux.scala 98:16]
  wire [4:0] _T_122 = _T_97 ? 5'h6 : _T_121; // @[Mux.scala 98:16]
  wire [4:0] _T_123 = _T_95 ? 5'h19 : _T_122; // @[Mux.scala 98:16]
  wire [4:0] _T_124 = _T_93 ? 5'h18 : _T_123; // @[Mux.scala 98:16]
  wire [4:0] _T_125 = _T_91 ? 5'h4 : _T_124; // @[Mux.scala 98:16]
  wire [4:0] _T_126 = _T_89 ? 5'h17 : _T_125; // @[Mux.scala 98:16]
  wire [4:0] _T_127 = _T_87 ? 5'h5 : _T_126; // @[Mux.scala 98:16]
  wire [4:0] _T_128 = _T_85 ? 5'hc : _T_127; // @[Mux.scala 98:16]
  wire [4:0] _T_129 = _T_83 ? 5'hf : _T_128; // @[Mux.scala 98:16]
  wire [4:0] _T_130 = _T_81 ? 5'he : _T_129; // @[Mux.scala 98:16]
  wire [4:0] _T_131 = _T_79 ? 5'h3 : _T_130; // @[Mux.scala 98:16]
  wire [4:0] _T_132 = _T_77 ? 5'h16 : _T_131; // @[Mux.scala 98:16]
  wire [4:0] _T_133 = _T_75 ? 5'h15 : _T_132; // @[Mux.scala 98:16]
  wire [4:0] _T_134 = _T_73 ? 5'h14 : _T_133; // @[Mux.scala 98:16]
  wire [4:0] _T_135 = _T_71 ? 5'h13 : _T_134; // @[Mux.scala 98:16]
  wire [4:0] _T_136 = _T_69 ? 5'h1 : _T_135; // @[Mux.scala 98:16]
  wire [4:0] _T_137 = _T_67 ? 5'h12 : _T_136; // @[Mux.scala 98:16]
  wire [4:0] _T_138 = _T_65 ? 5'h11 : _T_137; // @[Mux.scala 98:16]
  wire [4:0] _T_139 = _T_63 ? 5'h0 : _T_138; // @[Mux.scala 98:16]
  wire [4:0] _T_140 = _T_61 ? 5'h2 : _T_139; // @[Mux.scala 98:16]
  wire [4:0] _T_141 = _T_59 ? 5'h10 : _T_140; // @[Mux.scala 98:16]
  wire [4:0] _T_142 = _T_57 ? 5'hd : _T_141; // @[Mux.scala 98:16]
  wire [4:0] _T_143 = _T_55 ? 5'h7 : _T_142; // @[Mux.scala 98:16]
  wire [4:0] _T_144 = _T_53 ? 5'h3 : _T_143; // @[Mux.scala 98:16]
  wire [4:0] _T_145 = _T_51 ? 5'h0 : _T_144; // @[Mux.scala 98:16]
  wire [4:0] _T_146 = _T_49 ? 5'h0 : _T_145; // @[Mux.scala 98:16]
  wire [4:0] _T_147 = _T_47 ? 5'h0 : _T_146; // @[Mux.scala 98:16]
  wire [4:0] _T_148 = _T_17 ? 5'h0 : _T_147; // @[Mux.scala 98:16]
  wire [4:0] _T_149 = _T_43 ? 5'h0 : _T_148; // @[Mux.scala 98:16]
  wire [4:0] _T_150 = _T_41 ? 5'h0 : _T_149; // @[Mux.scala 98:16]
  wire [4:0] _T_151 = _T_39 ? 5'h9 : _T_150; // @[Mux.scala 98:16]
  wire [4:0] _T_152 = _T_37 ? 5'hf : _T_151; // @[Mux.scala 98:16]
  wire [4:0] _T_153 = _T_35 ? 5'he : _T_152; // @[Mux.scala 98:16]
  wire [4:0] _T_154 = _T_33 ? 5'h8 : _T_153; // @[Mux.scala 98:16]
  wire [4:0] _T_155 = _T_31 ? 5'hd : _T_154; // @[Mux.scala 98:16]
  wire [4:0] _T_156 = _T_29 ? 5'h4 : _T_155; // @[Mux.scala 98:16]
  wire [4:0] _T_157 = _T_27 ? 5'h2 : _T_156; // @[Mux.scala 98:16]
  wire [4:0] _T_158 = _T_25 ? 5'h6 : _T_157; // @[Mux.scala 98:16]
  wire [4:0] _T_159 = _T_23 ? 5'hc : _T_158; // @[Mux.scala 98:16]
  wire [4:0] _T_160 = _T_21 ? 5'h7 : _T_159; // @[Mux.scala 98:16]
  wire [4:0] _T_161 = _T_19 ? 5'h0 : _T_160; // @[Mux.scala 98:16]
  wire [4:0] _T_162 = _T_17 ? 5'h0 : _T_161; // @[Mux.scala 98:16]
  wire [4:0] _T_163 = _T_15 ? 5'h1f : _T_162; // @[Mux.scala 98:16]
  wire [4:0] _T_164 = _T_13 ? 5'h0 : _T_163; // @[Mux.scala 98:16]
  wire [4:0] _T_165 = _T_11 ? 5'ha : _T_164; // @[Mux.scala 98:16]
  wire [4:0] _T_166 = _T_9 ? 5'h0 : _T_165; // @[Mux.scala 98:16]
  wire [4:0] _T_167 = _T_7 ? 5'h0 : _T_166; // @[Mux.scala 98:16]
  wire [4:0] _T_168 = _T_5 ? 5'h0 : _T_167; // @[Mux.scala 98:16]
  wire [4:0] _T_169 = _T_3 ? 5'h0 : _T_168; // @[Mux.scala 98:16]
  assign io_ALUCtrl = _T_1 ? 5'h0 : _T_169; // @[ALUCtrl.scala 134:14]
endmodule
module ALUSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_AluSrc1,
  output [1:0]  io_AluSrc2
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[ALUSrcGen.scala 66:49]
  wire  _T_1 = 32'h2007033 == _T; // @[ALUSrcGen.scala 66:49]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[ALUSrcGen.scala 65:49]
  wire  _T_3 = 32'h1063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_5 = 32'h23 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_7 = 32'h6003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire [31:0] _T_8 = io_inst & 32'hfc00707f; // @[ALUSrcGen.scala 63:49]
  wire  _T_9 = 32'h1013 == _T_8; // @[ALUSrcGen.scala 63:49]
  wire  _T_11 = 32'h3033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_13 = 32'h200003b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_15 = 32'h5003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_17 = 32'h1b == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_19 = 32'h4000503b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_21 = 32'h3 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_23 = 32'h4033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_25 = 32'h5063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_27 = 32'h7033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_29 = 32'h200603b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_31 = 32'h2005033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_33 = 32'h2023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_35 = 32'h4003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_37 = 32'h2003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_39 = 32'h4000501b == _T; // @[ALUSrcGen.scala 63:49]
  wire  _T_41 = 32'h67 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_43 = 32'h4000003b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_45 = 32'h6063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_47 = 32'h3023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_49 = 32'h5013 == _T_8; // @[ALUSrcGen.scala 63:49]
  wire  _T_51 = 32'h1033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_53 = 32'h4063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_55 = 32'h101b == _T; // @[ALUSrcGen.scala 63:49]
  wire  _T_57 = 32'h200503b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_59 = 32'h3b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_61 = 32'h1023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_63 = 32'h4013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_65 = 32'h40000033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_67 = 32'h3013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_69 = 32'h2006033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_71 = 32'h1003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_73 = 32'h40005013 == _T_8; // @[ALUSrcGen.scala 63:49]
  wire  _T_75 = 32'h2000033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_77 = 32'h33 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_79 = 32'h3003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_81 = 32'h2033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_83 = 32'h200703b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_85 = 32'h5033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_87 = 32'h13 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_89 = 32'h501b == _T; // @[ALUSrcGen.scala 63:49]
  wire  _T_91 = 32'h103b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_93 = 32'h7063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_95 = 32'h6033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_97 = 32'h7013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_99 = 32'h503b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_101 = 32'h200403b == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_103 = 32'h2004033 == _T; // @[ALUSrcGen.scala 66:49]
  wire  _T_105 = 32'h63 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_107 = 32'h6013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire [31:0] _T_108 = io_inst & 32'h7f; // @[ALUSrcGen.scala 71:31]
  wire  _T_109 = 32'h17 == _T_108; // @[ALUSrcGen.scala 71:31]
  wire  _T_111 = 32'h37 == _T_108; // @[ALUSrcGen.scala 72:31]
  wire  _T_225 = _T_109 | _T_111; // @[Mux.scala 98:16]
  wire  _T_226 = _T_107 ? 1'h0 : _T_225; // @[Mux.scala 98:16]
  wire  _T_227 = _T_105 ? 1'h0 : _T_226; // @[Mux.scala 98:16]
  wire  _T_228 = _T_103 ? 1'h0 : _T_227; // @[Mux.scala 98:16]
  wire  _T_229 = _T_101 ? 1'h0 : _T_228; // @[Mux.scala 98:16]
  wire  _T_230 = _T_99 ? 1'h0 : _T_229; // @[Mux.scala 98:16]
  wire  _T_231 = _T_97 ? 1'h0 : _T_230; // @[Mux.scala 98:16]
  wire  _T_232 = _T_95 ? 1'h0 : _T_231; // @[Mux.scala 98:16]
  wire  _T_233 = _T_93 ? 1'h0 : _T_232; // @[Mux.scala 98:16]
  wire  _T_234 = _T_91 ? 1'h0 : _T_233; // @[Mux.scala 98:16]
  wire  _T_235 = _T_89 ? 1'h0 : _T_234; // @[Mux.scala 98:16]
  wire  _T_236 = _T_87 ? 1'h0 : _T_235; // @[Mux.scala 98:16]
  wire  _T_237 = _T_85 ? 1'h0 : _T_236; // @[Mux.scala 98:16]
  wire  _T_238 = _T_83 ? 1'h0 : _T_237; // @[Mux.scala 98:16]
  wire  _T_239 = _T_81 ? 1'h0 : _T_238; // @[Mux.scala 98:16]
  wire  _T_240 = _T_79 ? 1'h0 : _T_239; // @[Mux.scala 98:16]
  wire  _T_241 = _T_77 ? 1'h0 : _T_240; // @[Mux.scala 98:16]
  wire  _T_242 = _T_75 ? 1'h0 : _T_241; // @[Mux.scala 98:16]
  wire  _T_243 = _T_73 ? 1'h0 : _T_242; // @[Mux.scala 98:16]
  wire  _T_244 = _T_71 ? 1'h0 : _T_243; // @[Mux.scala 98:16]
  wire  _T_245 = _T_69 ? 1'h0 : _T_244; // @[Mux.scala 98:16]
  wire  _T_246 = _T_67 ? 1'h0 : _T_245; // @[Mux.scala 98:16]
  wire  _T_247 = _T_65 ? 1'h0 : _T_246; // @[Mux.scala 98:16]
  wire  _T_248 = _T_63 ? 1'h0 : _T_247; // @[Mux.scala 98:16]
  wire  _T_249 = _T_61 ? 1'h0 : _T_248; // @[Mux.scala 98:16]
  wire  _T_250 = _T_59 ? 1'h0 : _T_249; // @[Mux.scala 98:16]
  wire  _T_251 = _T_57 ? 1'h0 : _T_250; // @[Mux.scala 98:16]
  wire  _T_252 = _T_55 ? 1'h0 : _T_251; // @[Mux.scala 98:16]
  wire  _T_253 = _T_53 ? 1'h0 : _T_252; // @[Mux.scala 98:16]
  wire  _T_254 = _T_51 ? 1'h0 : _T_253; // @[Mux.scala 98:16]
  wire  _T_255 = _T_49 ? 1'h0 : _T_254; // @[Mux.scala 98:16]
  wire  _T_256 = _T_47 ? 1'h0 : _T_255; // @[Mux.scala 98:16]
  wire  _T_257 = _T_45 ? 1'h0 : _T_256; // @[Mux.scala 98:16]
  wire  _T_258 = _T_43 ? 1'h0 : _T_257; // @[Mux.scala 98:16]
  wire  _T_259 = _T_41 ? 1'h0 : _T_258; // @[Mux.scala 98:16]
  wire  _T_260 = _T_39 ? 1'h0 : _T_259; // @[Mux.scala 98:16]
  wire  _T_261 = _T_37 ? 1'h0 : _T_260; // @[Mux.scala 98:16]
  wire  _T_262 = _T_35 ? 1'h0 : _T_261; // @[Mux.scala 98:16]
  wire  _T_263 = _T_33 ? 1'h0 : _T_262; // @[Mux.scala 98:16]
  wire  _T_264 = _T_31 ? 1'h0 : _T_263; // @[Mux.scala 98:16]
  wire  _T_265 = _T_29 ? 1'h0 : _T_264; // @[Mux.scala 98:16]
  wire  _T_266 = _T_27 ? 1'h0 : _T_265; // @[Mux.scala 98:16]
  wire  _T_267 = _T_25 ? 1'h0 : _T_266; // @[Mux.scala 98:16]
  wire  _T_268 = _T_23 ? 1'h0 : _T_267; // @[Mux.scala 98:16]
  wire  _T_269 = _T_21 ? 1'h0 : _T_268; // @[Mux.scala 98:16]
  wire  _T_270 = _T_19 ? 1'h0 : _T_269; // @[Mux.scala 98:16]
  wire  _T_271 = _T_17 ? 1'h0 : _T_270; // @[Mux.scala 98:16]
  wire  _T_272 = _T_15 ? 1'h0 : _T_271; // @[Mux.scala 98:16]
  wire  _T_273 = _T_13 ? 1'h0 : _T_272; // @[Mux.scala 98:16]
  wire  _T_274 = _T_11 ? 1'h0 : _T_273; // @[Mux.scala 98:16]
  wire  _T_275 = _T_9 ? 1'h0 : _T_274; // @[Mux.scala 98:16]
  wire  _T_276 = _T_7 ? 1'h0 : _T_275; // @[Mux.scala 98:16]
  wire  _T_277 = _T_5 ? 1'h0 : _T_276; // @[Mux.scala 98:16]
  wire  _T_278 = _T_3 ? 1'h0 : _T_277; // @[Mux.scala 98:16]
  wire  _T_279 = _T_1 ? 1'h0 : _T_278; // @[Mux.scala 98:16]
  wire [1:0] _T_280 = _T_111 ? 2'h3 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_281 = _T_109 ? 2'h2 : _T_280; // @[Mux.scala 98:16]
  wire [1:0] _T_282 = _T_107 ? 2'h1 : _T_281; // @[Mux.scala 98:16]
  wire [1:0] _T_283 = _T_105 ? 2'h0 : _T_282; // @[Mux.scala 98:16]
  wire [1:0] _T_284 = _T_103 ? 2'h0 : _T_283; // @[Mux.scala 98:16]
  wire [1:0] _T_285 = _T_101 ? 2'h0 : _T_284; // @[Mux.scala 98:16]
  wire [1:0] _T_286 = _T_99 ? 2'h0 : _T_285; // @[Mux.scala 98:16]
  wire [1:0] _T_287 = _T_97 ? 2'h1 : _T_286; // @[Mux.scala 98:16]
  wire [1:0] _T_288 = _T_95 ? 2'h0 : _T_287; // @[Mux.scala 98:16]
  wire [1:0] _T_289 = _T_93 ? 2'h0 : _T_288; // @[Mux.scala 98:16]
  wire [1:0] _T_290 = _T_91 ? 2'h0 : _T_289; // @[Mux.scala 98:16]
  wire [1:0] _T_291 = _T_89 ? 2'h1 : _T_290; // @[Mux.scala 98:16]
  wire [1:0] _T_292 = _T_87 ? 2'h1 : _T_291; // @[Mux.scala 98:16]
  wire [1:0] _T_293 = _T_85 ? 2'h0 : _T_292; // @[Mux.scala 98:16]
  wire [1:0] _T_294 = _T_83 ? 2'h0 : _T_293; // @[Mux.scala 98:16]
  wire [1:0] _T_295 = _T_81 ? 2'h0 : _T_294; // @[Mux.scala 98:16]
  wire [1:0] _T_296 = _T_79 ? 2'h1 : _T_295; // @[Mux.scala 98:16]
  wire [1:0] _T_297 = _T_77 ? 2'h0 : _T_296; // @[Mux.scala 98:16]
  wire [1:0] _T_298 = _T_75 ? 2'h0 : _T_297; // @[Mux.scala 98:16]
  wire [1:0] _T_299 = _T_73 ? 2'h1 : _T_298; // @[Mux.scala 98:16]
  wire [1:0] _T_300 = _T_71 ? 2'h1 : _T_299; // @[Mux.scala 98:16]
  wire [1:0] _T_301 = _T_69 ? 2'h0 : _T_300; // @[Mux.scala 98:16]
  wire [1:0] _T_302 = _T_67 ? 2'h1 : _T_301; // @[Mux.scala 98:16]
  wire [1:0] _T_303 = _T_65 ? 2'h0 : _T_302; // @[Mux.scala 98:16]
  wire [1:0] _T_304 = _T_63 ? 2'h1 : _T_303; // @[Mux.scala 98:16]
  wire [1:0] _T_305 = _T_61 ? 2'h1 : _T_304; // @[Mux.scala 98:16]
  wire [1:0] _T_306 = _T_59 ? 2'h0 : _T_305; // @[Mux.scala 98:16]
  wire [1:0] _T_307 = _T_57 ? 2'h0 : _T_306; // @[Mux.scala 98:16]
  wire [1:0] _T_308 = _T_55 ? 2'h1 : _T_307; // @[Mux.scala 98:16]
  wire [1:0] _T_309 = _T_53 ? 2'h0 : _T_308; // @[Mux.scala 98:16]
  wire [1:0] _T_310 = _T_51 ? 2'h0 : _T_309; // @[Mux.scala 98:16]
  wire [1:0] _T_311 = _T_49 ? 2'h1 : _T_310; // @[Mux.scala 98:16]
  wire [1:0] _T_312 = _T_47 ? 2'h1 : _T_311; // @[Mux.scala 98:16]
  wire [1:0] _T_313 = _T_45 ? 2'h0 : _T_312; // @[Mux.scala 98:16]
  wire [1:0] _T_314 = _T_43 ? 2'h0 : _T_313; // @[Mux.scala 98:16]
  wire [1:0] _T_315 = _T_41 ? 2'h1 : _T_314; // @[Mux.scala 98:16]
  wire [1:0] _T_316 = _T_39 ? 2'h1 : _T_315; // @[Mux.scala 98:16]
  wire [1:0] _T_317 = _T_37 ? 2'h1 : _T_316; // @[Mux.scala 98:16]
  wire [1:0] _T_318 = _T_35 ? 2'h1 : _T_317; // @[Mux.scala 98:16]
  wire [1:0] _T_319 = _T_33 ? 2'h1 : _T_318; // @[Mux.scala 98:16]
  wire [1:0] _T_320 = _T_31 ? 2'h0 : _T_319; // @[Mux.scala 98:16]
  wire [1:0] _T_321 = _T_29 ? 2'h0 : _T_320; // @[Mux.scala 98:16]
  wire [1:0] _T_322 = _T_27 ? 2'h0 : _T_321; // @[Mux.scala 98:16]
  wire [1:0] _T_323 = _T_25 ? 2'h0 : _T_322; // @[Mux.scala 98:16]
  wire [1:0] _T_324 = _T_23 ? 2'h0 : _T_323; // @[Mux.scala 98:16]
  wire [1:0] _T_325 = _T_21 ? 2'h1 : _T_324; // @[Mux.scala 98:16]
  wire [1:0] _T_326 = _T_19 ? 2'h0 : _T_325; // @[Mux.scala 98:16]
  wire [1:0] _T_327 = _T_17 ? 2'h1 : _T_326; // @[Mux.scala 98:16]
  wire [1:0] _T_328 = _T_15 ? 2'h1 : _T_327; // @[Mux.scala 98:16]
  wire [1:0] _T_329 = _T_13 ? 2'h0 : _T_328; // @[Mux.scala 98:16]
  wire [1:0] _T_330 = _T_11 ? 2'h0 : _T_329; // @[Mux.scala 98:16]
  wire [1:0] _T_331 = _T_9 ? 2'h1 : _T_330; // @[Mux.scala 98:16]
  wire [1:0] _T_332 = _T_7 ? 2'h1 : _T_331; // @[Mux.scala 98:16]
  wire [1:0] _T_333 = _T_5 ? 2'h1 : _T_332; // @[Mux.scala 98:16]
  wire [1:0] _T_334 = _T_3 ? 2'h0 : _T_333; // @[Mux.scala 98:16]
  assign io_AluSrc1 = {{1'd0}, _T_279}; // @[ALUSrcGen.scala 90:14]
  assign io_AluSrc2 = _T_1 ? 2'h0 : _T_334; // @[ALUSrcGen.scala 91:14]
endmodule
module memWriteMGen(
  input  [31:0] io_inst,
  output        io_memWriteM
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memWriteMGen.scala 19:49]
  wire  _T_1 = 32'h23 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_3 = 32'h2023 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_5 = 32'h3023 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_7 = 32'h1023 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_9 = _T_5 | _T_7; // @[Mux.scala 98:16]
  wire  _T_10 = _T_3 | _T_9; // @[Mux.scala 98:16]
  assign io_memWriteM = _T_1 | _T_10; // @[memWriteMGen.scala 25:16]
endmodule
module memWriteMaskGen(
  input  [31:0] io_inst,
  output [7:0]  io_mask
);
  wire  _T_1 = 3'h0 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_2 = _T_1 ? 8'h1 : 8'h0; // @[Mux.scala 80:57]
  wire  _T_3 = 3'h1 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_4 = _T_3 ? 8'h3 : _T_2; // @[Mux.scala 80:57]
  wire  _T_5 = 3'h2 == io_inst[14:12]; // @[Mux.scala 80:60]
  wire [7:0] _T_6 = _T_5 ? 8'hf : _T_4; // @[Mux.scala 80:57]
  wire  _T_7 = 3'h3 == io_inst[14:12]; // @[Mux.scala 80:60]
  assign io_mask = _T_7 ? 8'hff : _T_6; // @[memWriteMaskGen.scala 19:11]
endmodule
module memReadNumGen(
  input  [31:0] io_inst,
  output [2:0]  io_memReadNum
);
  assign io_memReadNum = io_inst[14:12]; // @[memReadNumGen.scala 22:17]
endmodule
module dnpcSrcGen(
  input  [31:0] io_inst,
  output        io_dnpcSrc
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 25:49]
  wire  _T_1 = 32'h1063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_3 = 32'h5063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_5 = 32'h6063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_7 = 32'h4063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_9 = 32'h7063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_11 = 32'h63 == _T; // @[npcSrcGen.scala 25:49]
  wire [31:0] _T_12 = io_inst & 32'h7f; // @[npcSrcGen.scala 30:31]
  wire  _T_13 = 32'h6f == _T_12; // @[npcSrcGen.scala 30:31]
  wire  _T_18 = _T_11 | _T_13; // @[Mux.scala 98:16]
  wire  _T_19 = _T_9 | _T_18; // @[Mux.scala 98:16]
  wire  _T_20 = _T_7 | _T_19; // @[Mux.scala 98:16]
  wire  _T_21 = _T_5 | _T_20; // @[Mux.scala 98:16]
  wire  _T_22 = _T_3 | _T_21; // @[Mux.scala 98:16]
  assign io_dnpcSrc = _T_1 | _T_22; // @[npcSrcGen.scala 33:14]
endmodule
module jumpGen(
  input  [31:0] io_inst,
  output        io_jump
);
  wire [31:0] _T = io_inst & 32'h7f; // @[npcSrcGen.scala 46:14]
  wire  _T_1 = 32'h6f == _T; // @[npcSrcGen.scala 46:14]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[npcSrcGen.scala 47:14]
  wire  _T_3 = 32'h67 == _T_2; // @[npcSrcGen.scala 47:14]
  assign io_jump = _T_1 | _T_3; // @[npcSrcGen.scala 50:11]
endmodule
module branchGen(
  input  [31:0] io_inst,
  output        io_branch
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 66:47]
  wire  _T_1 = 32'h1063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_3 = 32'h5063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_5 = 32'h6063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_7 = 32'h4063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_9 = 32'h7063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_11 = 32'h63 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_13 = _T_9 | _T_11; // @[Mux.scala 98:16]
  wire  _T_14 = _T_7 | _T_13; // @[Mux.scala 98:16]
  wire  _T_15 = _T_5 | _T_14; // @[Mux.scala 98:16]
  wire  _T_16 = _T_3 | _T_15; // @[Mux.scala 98:16]
  assign io_branch = _T_1 | _T_16; // @[npcSrcGen.scala 72:13]
endmodule
module regEnGen(
  input  [31:0] io_inst,
  output        io_regEn
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[regEnGen.scala 35:45]
  wire  _T_1 = 32'h2007033 == _T; // @[regEnGen.scala 35:45]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[regEnGen.scala 37:45]
  wire  _T_3 = 32'h1063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_5 = 32'h23 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_7 = 32'h6003 == _T_2; // @[regEnGen.scala 33:45]
  wire [31:0] _T_8 = io_inst & 32'hfc00707f; // @[regEnGen.scala 33:45]
  wire  _T_9 = 32'h1013 == _T_8; // @[regEnGen.scala 33:45]
  wire  _T_11 = 32'h3033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_13 = 32'h200003b == _T; // @[regEnGen.scala 35:45]
  wire  _T_15 = 32'h5003 == _T_2; // @[regEnGen.scala 33:45]
  wire [31:0] _T_16 = io_inst & 32'h7f; // @[regEnGen.scala 32:45]
  wire  _T_17 = 32'h17 == _T_16; // @[regEnGen.scala 32:45]
  wire  _T_19 = 32'h1b == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_21 = 32'h4000503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_23 = 32'h3 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_25 = 32'h4033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_27 = 32'h5063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_29 = 32'h7033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_31 = 32'h200603b == _T; // @[regEnGen.scala 35:45]
  wire  _T_33 = 32'h2005033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_35 = 32'h2023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_37 = 32'h4003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_39 = 32'h2003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_41 = 32'h6f == _T_16; // @[regEnGen.scala 34:45]
  wire  _T_43 = 32'h4000501b == _T; // @[regEnGen.scala 33:45]
  wire  _T_45 = 32'h67 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_47 = 32'h4000003b == _T; // @[regEnGen.scala 35:45]
  wire  _T_49 = 32'h6063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_51 = 32'h3023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_53 = 32'h5013 == _T_8; // @[regEnGen.scala 33:45]
  wire  _T_55 = 32'h1033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_57 = 32'h4063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_59 = 32'h101b == _T; // @[regEnGen.scala 33:45]
  wire  _T_61 = 32'h200503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_63 = 32'h3b == _T; // @[regEnGen.scala 35:45]
  wire  _T_65 = 32'h37 == _T_16; // @[regEnGen.scala 32:45]
  wire  _T_67 = 32'h1023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_69 = 32'h4013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_71 = 32'h40000033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_73 = 32'h3013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_75 = 32'h2006033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_77 = 32'h1003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_79 = 32'h40005013 == _T_8; // @[regEnGen.scala 33:45]
  wire  _T_81 = 32'h2000033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_83 = 32'h33 == _T; // @[regEnGen.scala 35:45]
  wire  _T_85 = 32'h3003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_87 = 32'h2033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_89 = 32'h200703b == _T; // @[regEnGen.scala 35:45]
  wire  _T_91 = 32'h5033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_93 = 32'h13 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_95 = 32'h501b == _T; // @[regEnGen.scala 33:45]
  wire  _T_97 = 32'h103b == _T; // @[regEnGen.scala 35:45]
  wire  _T_99 = 32'h7063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_101 = 32'h6033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_103 = 32'h7013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_105 = 32'h503b == _T; // @[regEnGen.scala 35:45]
  wire  _T_107 = 32'h200403b == _T; // @[regEnGen.scala 35:45]
  wire  _T_109 = 32'h2004033 == _T; // @[regEnGen.scala 35:45]
  wire  _T_111 = 32'h63 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_113 = 32'h6013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_115 = _T_111 ? 1'h0 : _T_113; // @[Mux.scala 98:16]
  wire  _T_116 = _T_109 | _T_115; // @[Mux.scala 98:16]
  wire  _T_117 = _T_107 | _T_116; // @[Mux.scala 98:16]
  wire  _T_118 = _T_105 | _T_117; // @[Mux.scala 98:16]
  wire  _T_119 = _T_103 | _T_118; // @[Mux.scala 98:16]
  wire  _T_120 = _T_101 | _T_119; // @[Mux.scala 98:16]
  wire  _T_121 = _T_99 ? 1'h0 : _T_120; // @[Mux.scala 98:16]
  wire  _T_122 = _T_97 | _T_121; // @[Mux.scala 98:16]
  wire  _T_123 = _T_95 | _T_122; // @[Mux.scala 98:16]
  wire  _T_124 = _T_93 | _T_123; // @[Mux.scala 98:16]
  wire  _T_125 = _T_91 | _T_124; // @[Mux.scala 98:16]
  wire  _T_126 = _T_89 | _T_125; // @[Mux.scala 98:16]
  wire  _T_127 = _T_87 | _T_126; // @[Mux.scala 98:16]
  wire  _T_128 = _T_85 | _T_127; // @[Mux.scala 98:16]
  wire  _T_129 = _T_83 | _T_128; // @[Mux.scala 98:16]
  wire  _T_130 = _T_81 | _T_129; // @[Mux.scala 98:16]
  wire  _T_131 = _T_79 | _T_130; // @[Mux.scala 98:16]
  wire  _T_132 = _T_77 | _T_131; // @[Mux.scala 98:16]
  wire  _T_133 = _T_75 | _T_132; // @[Mux.scala 98:16]
  wire  _T_134 = _T_73 | _T_133; // @[Mux.scala 98:16]
  wire  _T_135 = _T_71 | _T_134; // @[Mux.scala 98:16]
  wire  _T_136 = _T_69 | _T_135; // @[Mux.scala 98:16]
  wire  _T_137 = _T_67 ? 1'h0 : _T_136; // @[Mux.scala 98:16]
  wire  _T_138 = _T_65 | _T_137; // @[Mux.scala 98:16]
  wire  _T_139 = _T_63 | _T_138; // @[Mux.scala 98:16]
  wire  _T_140 = _T_61 | _T_139; // @[Mux.scala 98:16]
  wire  _T_141 = _T_59 | _T_140; // @[Mux.scala 98:16]
  wire  _T_142 = _T_57 ? 1'h0 : _T_141; // @[Mux.scala 98:16]
  wire  _T_143 = _T_55 | _T_142; // @[Mux.scala 98:16]
  wire  _T_144 = _T_53 | _T_143; // @[Mux.scala 98:16]
  wire  _T_145 = _T_51 ? 1'h0 : _T_144; // @[Mux.scala 98:16]
  wire  _T_146 = _T_49 ? 1'h0 : _T_145; // @[Mux.scala 98:16]
  wire  _T_147 = _T_47 | _T_146; // @[Mux.scala 98:16]
  wire  _T_148 = _T_45 | _T_147; // @[Mux.scala 98:16]
  wire  _T_149 = _T_43 | _T_148; // @[Mux.scala 98:16]
  wire  _T_150 = _T_41 | _T_149; // @[Mux.scala 98:16]
  wire  _T_151 = _T_39 | _T_150; // @[Mux.scala 98:16]
  wire  _T_152 = _T_37 | _T_151; // @[Mux.scala 98:16]
  wire  _T_153 = _T_35 ? 1'h0 : _T_152; // @[Mux.scala 98:16]
  wire  _T_154 = _T_33 | _T_153; // @[Mux.scala 98:16]
  wire  _T_155 = _T_31 | _T_154; // @[Mux.scala 98:16]
  wire  _T_156 = _T_29 | _T_155; // @[Mux.scala 98:16]
  wire  _T_157 = _T_27 ? 1'h0 : _T_156; // @[Mux.scala 98:16]
  wire  _T_158 = _T_25 | _T_157; // @[Mux.scala 98:16]
  wire  _T_159 = _T_23 | _T_158; // @[Mux.scala 98:16]
  wire  _T_160 = _T_21 | _T_159; // @[Mux.scala 98:16]
  wire  _T_161 = _T_19 | _T_160; // @[Mux.scala 98:16]
  wire  _T_162 = _T_17 | _T_161; // @[Mux.scala 98:16]
  wire  _T_163 = _T_15 | _T_162; // @[Mux.scala 98:16]
  wire  _T_164 = _T_13 | _T_163; // @[Mux.scala 98:16]
  wire  _T_165 = _T_11 | _T_164; // @[Mux.scala 98:16]
  wire  _T_166 = _T_9 | _T_165; // @[Mux.scala 98:16]
  wire  _T_167 = _T_7 | _T_166; // @[Mux.scala 98:16]
  wire  _T_168 = _T_5 ? 1'h0 : _T_167; // @[Mux.scala 98:16]
  wire  _T_169 = _T_3 ? 1'h0 : _T_168; // @[Mux.scala 98:16]
  assign io_regEn = _T_1 | _T_169; // @[regEnGen.scala 43:12]
endmodule
module ResultSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_ResultSrc
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[ResultSrcGen.scala 39:44]
  wire  _T_1 = 32'h2007033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_3 = 32'h3033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_5 = 32'h200003b == _T; // @[ResultSrcGen.scala 39:44]
  wire [31:0] _T_6 = io_inst & 32'h7f; // @[ResultSrcGen.scala 37:44]
  wire  _T_7 = 32'h17 == _T_6; // @[ResultSrcGen.scala 37:44]
  wire  _T_9 = 32'h4000503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_11 = 32'h4033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_13 = 32'h7033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_15 = 32'h200603b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_17 = 32'h2005033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_19 = 32'h6f == _T_6; // @[ResultSrcGen.scala 38:44]
  wire  _T_21 = 32'h4000003b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_23 = 32'h1033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_25 = 32'h200503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_27 = 32'h3b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_29 = 32'h37 == _T_6; // @[ResultSrcGen.scala 37:44]
  wire  _T_31 = 32'h40000033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_33 = 32'h2006033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_35 = 32'h2000033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_37 = 32'h33 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_39 = 32'h2033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_41 = 32'h200703b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_43 = 32'h5033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_45 = 32'h103b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_47 = 32'h6033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_49 = 32'h503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_51 = 32'h200403b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_53 = 32'h2004033 == _T; // @[ResultSrcGen.scala 39:44]
  wire [31:0] _T_54 = io_inst & 32'h707f; // @[ResultSrcGen.scala 44:26]
  wire  _T_55 = 32'h13 == _T_54; // @[ResultSrcGen.scala 44:26]
  wire  _T_57 = 32'h67 == _T_54; // @[ResultSrcGen.scala 45:26]
  wire  _T_61 = 32'h3003 == _T_54; // @[ResultSrcGen.scala 47:26]
  wire  _T_63 = 32'h4003 == _T_54; // @[ResultSrcGen.scala 48:26]
  wire  _T_65 = 32'h3013 == _T_54; // @[ResultSrcGen.scala 49:26]
  wire  _T_67 = 32'h501b == _T; // @[ResultSrcGen.scala 50:26]
  wire [31:0] _T_68 = io_inst & 32'hfc00707f; // @[ResultSrcGen.scala 51:26]
  wire  _T_69 = 32'h1013 == _T_68; // @[ResultSrcGen.scala 51:26]
  wire  _T_71 = 32'h7013 == _T_54; // @[ResultSrcGen.scala 52:26]
  wire  _T_73 = 32'h4013 == _T_54; // @[ResultSrcGen.scala 53:26]
  wire  _T_75 = 32'h1b == _T_54; // @[ResultSrcGen.scala 54:26]
  wire  _T_77 = 32'h5013 == _T_68; // @[ResultSrcGen.scala 55:26]
  wire  _T_79 = 32'h101b == _T; // @[ResultSrcGen.scala 56:26]
  wire  _T_81 = 32'h4000501b == _T; // @[ResultSrcGen.scala 57:26]
  wire  _T_83 = 32'h40005013 == _T_68; // @[ResultSrcGen.scala 58:26]
  wire  _T_85 = 32'h6013 == _T_54; // @[ResultSrcGen.scala 59:26]
  wire  _T_87 = 32'h1003 == _T_54; // @[ResultSrcGen.scala 60:26]
  wire  _T_89 = 32'h2003 == _T_54; // @[ResultSrcGen.scala 61:26]
  wire  _T_91 = 32'h5003 == _T_54; // @[ResultSrcGen.scala 62:26]
  wire  _T_93 = 32'h6003 == _T_54; // @[ResultSrcGen.scala 63:26]
  wire  _T_95 = 32'h3 == _T_54; // @[ResultSrcGen.scala 64:26]
  wire [1:0] _T_102 = _T_95 ? 2'h2 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_103 = _T_93 ? 2'h2 : _T_102; // @[Mux.scala 98:16]
  wire [1:0] _T_104 = _T_91 ? 2'h2 : _T_103; // @[Mux.scala 98:16]
  wire [1:0] _T_105 = _T_89 ? 2'h2 : _T_104; // @[Mux.scala 98:16]
  wire [1:0] _T_106 = _T_87 ? 2'h2 : _T_105; // @[Mux.scala 98:16]
  wire [1:0] _T_107 = _T_85 ? 2'h0 : _T_106; // @[Mux.scala 98:16]
  wire [1:0] _T_108 = _T_83 ? 2'h0 : _T_107; // @[Mux.scala 98:16]
  wire [1:0] _T_109 = _T_81 ? 2'h0 : _T_108; // @[Mux.scala 98:16]
  wire [1:0] _T_110 = _T_79 ? 2'h0 : _T_109; // @[Mux.scala 98:16]
  wire [1:0] _T_111 = _T_77 ? 2'h0 : _T_110; // @[Mux.scala 98:16]
  wire [1:0] _T_112 = _T_75 ? 2'h0 : _T_111; // @[Mux.scala 98:16]
  wire [1:0] _T_113 = _T_73 ? 2'h0 : _T_112; // @[Mux.scala 98:16]
  wire [1:0] _T_114 = _T_71 ? 2'h0 : _T_113; // @[Mux.scala 98:16]
  wire [1:0] _T_115 = _T_69 ? 2'h0 : _T_114; // @[Mux.scala 98:16]
  wire [1:0] _T_116 = _T_67 ? 2'h0 : _T_115; // @[Mux.scala 98:16]
  wire [1:0] _T_117 = _T_65 ? 2'h0 : _T_116; // @[Mux.scala 98:16]
  wire [1:0] _T_118 = _T_63 ? 2'h2 : _T_117; // @[Mux.scala 98:16]
  wire [1:0] _T_119 = _T_61 ? 2'h2 : _T_118; // @[Mux.scala 98:16]
  wire [1:0] _T_120 = _T_57 ? 2'h1 : _T_119; // @[Mux.scala 98:16]
  wire [1:0] _T_121 = _T_57 ? 2'h1 : _T_120; // @[Mux.scala 98:16]
  wire [1:0] _T_122 = _T_55 ? 2'h0 : _T_121; // @[Mux.scala 98:16]
  wire [1:0] _T_123 = _T_53 ? 2'h0 : _T_122; // @[Mux.scala 98:16]
  wire [1:0] _T_124 = _T_51 ? 2'h0 : _T_123; // @[Mux.scala 98:16]
  wire [1:0] _T_125 = _T_49 ? 2'h0 : _T_124; // @[Mux.scala 98:16]
  wire [1:0] _T_126 = _T_47 ? 2'h0 : _T_125; // @[Mux.scala 98:16]
  wire [1:0] _T_127 = _T_45 ? 2'h0 : _T_126; // @[Mux.scala 98:16]
  wire [1:0] _T_128 = _T_43 ? 2'h0 : _T_127; // @[Mux.scala 98:16]
  wire [1:0] _T_129 = _T_41 ? 2'h0 : _T_128; // @[Mux.scala 98:16]
  wire [1:0] _T_130 = _T_39 ? 2'h0 : _T_129; // @[Mux.scala 98:16]
  wire [1:0] _T_131 = _T_37 ? 2'h0 : _T_130; // @[Mux.scala 98:16]
  wire [1:0] _T_132 = _T_35 ? 2'h0 : _T_131; // @[Mux.scala 98:16]
  wire [1:0] _T_133 = _T_33 ? 2'h0 : _T_132; // @[Mux.scala 98:16]
  wire [1:0] _T_134 = _T_31 ? 2'h0 : _T_133; // @[Mux.scala 98:16]
  wire [1:0] _T_135 = _T_29 ? 2'h0 : _T_134; // @[Mux.scala 98:16]
  wire [1:0] _T_136 = _T_27 ? 2'h0 : _T_135; // @[Mux.scala 98:16]
  wire [1:0] _T_137 = _T_25 ? 2'h0 : _T_136; // @[Mux.scala 98:16]
  wire [1:0] _T_138 = _T_23 ? 2'h0 : _T_137; // @[Mux.scala 98:16]
  wire [1:0] _T_139 = _T_21 ? 2'h0 : _T_138; // @[Mux.scala 98:16]
  wire [1:0] _T_140 = _T_19 ? 2'h1 : _T_139; // @[Mux.scala 98:16]
  wire [1:0] _T_141 = _T_17 ? 2'h0 : _T_140; // @[Mux.scala 98:16]
  wire [1:0] _T_142 = _T_15 ? 2'h0 : _T_141; // @[Mux.scala 98:16]
  wire [1:0] _T_143 = _T_13 ? 2'h0 : _T_142; // @[Mux.scala 98:16]
  wire [1:0] _T_144 = _T_11 ? 2'h0 : _T_143; // @[Mux.scala 98:16]
  wire [1:0] _T_145 = _T_9 ? 2'h0 : _T_144; // @[Mux.scala 98:16]
  wire [1:0] _T_146 = _T_7 ? 2'h0 : _T_145; // @[Mux.scala 98:16]
  wire [1:0] _T_147 = _T_5 ? 2'h0 : _T_146; // @[Mux.scala 98:16]
  wire [1:0] _T_148 = _T_3 ? 2'h0 : _T_147; // @[Mux.scala 98:16]
  assign io_ResultSrc = _T_1 ? 2'h0 : _T_148; // @[ResultSrcGen.scala 68:16]
endmodule
module CtrlUnit(
  input  [31:0] io_inst,
  output [1:0]  io_CtrlS_AluSrc1,
  output [1:0]  io_CtrlS_AluSrc2,
  output [4:0]  io_CtrlS_ALUCtrl,
  output        io_CtrlS_memWriteM,
  output [7:0]  io_CtrlS_memWriteMask,
  output [2:0]  io_CtrlS_memReadNum,
  output        io_CtrlS_dnpcSrc,
  output        io_CtrlS_jump,
  output        io_CtrlS_branch,
  output        io_CtrlS_regEn,
  output [1:0]  io_CtrlS_ResultSrc,
  output        io_CtrlS_fencei
);
  wire [31:0] ALUCtrl_ins_io_inst; // @[CtrlUnit.scala 33:26]
  wire [4:0] ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 33:26]
  wire [31:0] ALUSrcGen_ins_io_inst; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 37:29]
  wire [31:0] memWriteMGen_ins_io_inst; // @[CtrlUnit.scala 42:32]
  wire  memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 42:32]
  wire [31:0] memWriteMaskGen_ins_io_inst; // @[CtrlUnit.scala 46:35]
  wire [7:0] memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 46:35]
  wire [31:0] memReadNumGen_ins_io_inst; // @[CtrlUnit.scala 50:33]
  wire [2:0] memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 50:33]
  wire [31:0] dnpcSrcGen_ins_io_inst; // @[CtrlUnit.scala 54:32]
  wire  dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 54:32]
  wire [31:0] jumpGen_ins_io_inst; // @[CtrlUnit.scala 58:27]
  wire  jumpGen_ins_io_jump; // @[CtrlUnit.scala 58:27]
  wire [31:0] branchGen_ins_io_inst; // @[CtrlUnit.scala 62:29]
  wire  branchGen_ins_io_branch; // @[CtrlUnit.scala 62:29]
  wire [31:0] regEnGen_ins_io_inst; // @[CtrlUnit.scala 67:28]
  wire  regEnGen_ins_io_regEn; // @[CtrlUnit.scala 67:28]
  wire [31:0] ResultSrcGen_ins_io_inst; // @[CtrlUnit.scala 71:32]
  wire [1:0] ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 71:32]
  wire [31:0] _T = io_inst & 32'h707f; // @[CtrlUnit.scala 75:30]
  ALUCtrl ALUCtrl_ins ( // @[CtrlUnit.scala 33:26]
    .io_inst(ALUCtrl_ins_io_inst),
    .io_ALUCtrl(ALUCtrl_ins_io_ALUCtrl)
  );
  ALUSrcGen ALUSrcGen_ins ( // @[CtrlUnit.scala 37:29]
    .io_inst(ALUSrcGen_ins_io_inst),
    .io_AluSrc1(ALUSrcGen_ins_io_AluSrc1),
    .io_AluSrc2(ALUSrcGen_ins_io_AluSrc2)
  );
  memWriteMGen memWriteMGen_ins ( // @[CtrlUnit.scala 42:32]
    .io_inst(memWriteMGen_ins_io_inst),
    .io_memWriteM(memWriteMGen_ins_io_memWriteM)
  );
  memWriteMaskGen memWriteMaskGen_ins ( // @[CtrlUnit.scala 46:35]
    .io_inst(memWriteMaskGen_ins_io_inst),
    .io_mask(memWriteMaskGen_ins_io_mask)
  );
  memReadNumGen memReadNumGen_ins ( // @[CtrlUnit.scala 50:33]
    .io_inst(memReadNumGen_ins_io_inst),
    .io_memReadNum(memReadNumGen_ins_io_memReadNum)
  );
  dnpcSrcGen dnpcSrcGen_ins ( // @[CtrlUnit.scala 54:32]
    .io_inst(dnpcSrcGen_ins_io_inst),
    .io_dnpcSrc(dnpcSrcGen_ins_io_dnpcSrc)
  );
  jumpGen jumpGen_ins ( // @[CtrlUnit.scala 58:27]
    .io_inst(jumpGen_ins_io_inst),
    .io_jump(jumpGen_ins_io_jump)
  );
  branchGen branchGen_ins ( // @[CtrlUnit.scala 62:29]
    .io_inst(branchGen_ins_io_inst),
    .io_branch(branchGen_ins_io_branch)
  );
  regEnGen regEnGen_ins ( // @[CtrlUnit.scala 67:28]
    .io_inst(regEnGen_ins_io_inst),
    .io_regEn(regEnGen_ins_io_regEn)
  );
  ResultSrcGen ResultSrcGen_ins ( // @[CtrlUnit.scala 71:32]
    .io_inst(ResultSrcGen_ins_io_inst),
    .io_ResultSrc(ResultSrcGen_ins_io_ResultSrc)
  );
  assign io_CtrlS_AluSrc1 = ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 39:20]
  assign io_CtrlS_AluSrc2 = ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 40:20]
  assign io_CtrlS_ALUCtrl = ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 35:20]
  assign io_CtrlS_memWriteM = memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 44:22]
  assign io_CtrlS_memWriteMask = memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 48:25]
  assign io_CtrlS_memReadNum = memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 52:23]
  assign io_CtrlS_dnpcSrc = dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 56:20]
  assign io_CtrlS_jump = jumpGen_ins_io_jump; // @[CtrlUnit.scala 60:17]
  assign io_CtrlS_branch = branchGen_ins_io_branch; // @[CtrlUnit.scala 64:19]
  assign io_CtrlS_regEn = regEnGen_ins_io_regEn; // @[CtrlUnit.scala 69:18]
  assign io_CtrlS_ResultSrc = ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 73:22]
  assign io_CtrlS_fencei = 32'h100f == _T; // @[CtrlUnit.scala 75:19]
  assign ALUCtrl_ins_io_inst = io_inst; // @[CtrlUnit.scala 34:23]
  assign ALUSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 38:25]
  assign memWriteMGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 43:28]
  assign memWriteMaskGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 47:31]
  assign memReadNumGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 51:29]
  assign dnpcSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 55:26]
  assign jumpGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 59:23]
  assign branchGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 63:25]
  assign regEnGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 68:24]
  assign ResultSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 72:28]
endmodule
module csrCtrl(
  input  [31:0] io_inst,
  output        io_CSRCtrlIf_csrrwen,
  output        io_CSRCtrlIf_csrswen,
  output        io_CSRCtrlIf_csrrsien,
  output        io_CSRCtrlIf_csrrcien,
  output        io_CSRCtrlIf_csrrcen,
  output        io_CSRCtrlIf_csrrwien,
  output        io_CSRCtrlIf_ecall,
  output        io_CSRCtrlIf_rfen,
  output        io_CSRCtrlIf_mepc2pc
);
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[csrCtrl.scala 43:35]
  wire  _T_3 = 32'h1073 == _T_2; // @[csrCtrl.scala 43:35]
  wire  _T_5 = 32'h2073 == _T_2; // @[csrCtrl.scala 44:35]
  wire  _T_7 = 32'h6073 == _T_2; // @[csrCtrl.scala 45:36]
  wire  _T_9 = 32'h7073 == _T_2; // @[csrCtrl.scala 46:36]
  wire  _T_11 = 32'h3073 == _T_2; // @[csrCtrl.scala 47:35]
  wire  _T_18 = _T_3 | _T_5; // @[csrCtrl.scala 50:41]
  wire  _T_21 = _T_18 | _T_7; // @[csrCtrl.scala 50:61]
  wire  _T_24 = _T_21 | _T_9; // @[csrCtrl.scala 50:81]
  assign io_CSRCtrlIf_csrrwen = 32'h1073 == _T_2; // @[csrCtrl.scala 43:24]
  assign io_CSRCtrlIf_csrswen = 32'h2073 == _T_2; // @[csrCtrl.scala 44:24]
  assign io_CSRCtrlIf_csrrsien = 32'h6073 == _T_2; // @[csrCtrl.scala 45:25]
  assign io_CSRCtrlIf_csrrcien = 32'h7073 == _T_2; // @[csrCtrl.scala 46:25]
  assign io_CSRCtrlIf_csrrcen = 32'h3073 == _T_2; // @[csrCtrl.scala 47:24]
  assign io_CSRCtrlIf_csrrwien = 32'h5073 == _T_2; // @[csrCtrl.scala 48:25]
  assign io_CSRCtrlIf_ecall = 32'h73 == io_inst; // @[csrCtrl.scala 40:22]
  assign io_CSRCtrlIf_rfen = _T_24 | _T_11; // @[csrCtrl.scala 50:21]
  assign io_CSRCtrlIf_mepc2pc = 32'h30200073 == io_inst; // @[csrCtrl.scala 52:24]
endmodule
module riscv(
  input         clock,
  input         reset,
  output        io_instIO_valid,
  input         io_instIO_ready,
  input  [63:0] io_instIO_data_read,
  output [31:0] io_instIO_addr,
  output        io_dataIO_valid,
  input         io_dataIO_ready,
  input  [63:0] io_dataIO_data_read,
  output [63:0] io_dataIO_data_write,
  output        io_dataIO_wen,
  output [31:0] io_dataIO_addr,
  output [1:0]  io_dataIO_rsize,
  output [7:0]  io_dataIO_mask,
  input         intrTimeCnt_0,
  output        startTimeCnt,
  output        block2_0,
  output        fencei_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [383:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [191:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[riscv.scala 31:19]
  wire  ifu_reset; // @[riscv.scala 31:19]
  wire [31:0] ifu_io_instIn; // @[riscv.scala 31:19]
  wire [31:0] ifu_io_instOut; // @[riscv.scala 31:19]
  wire [31:0] ifu_io_pc; // @[riscv.scala 31:19]
  wire [31:0] ifu_io_snpc; // @[riscv.scala 31:19]
  wire [31:0] ifu_io_dnpc; // @[riscv.scala 31:19]
  wire  ifu_io_jump; // @[riscv.scala 31:19]
  wire  ifu_intrTimeCnt_0; // @[riscv.scala 31:19]
  wire  ifu_hazardPCBlock_0; // @[riscv.scala 31:19]
  wire  ifu_block1_0; // @[riscv.scala 31:19]
  wire  ifu_block23_0; // @[riscv.scala 31:19]
  wire  idu_clock; // @[riscv.scala 32:19]
  wire [31:0] idu_io_pc; // @[riscv.scala 32:19]
  wire [31:0] idu_io_inst; // @[riscv.scala 32:19]
  wire  idu_io_regEn; // @[riscv.scala 32:19]
  wire [63:0] idu_io_dataEx_imme; // @[riscv.scala 32:19]
  wire [63:0] idu_io_dataEx_dOut1; // @[riscv.scala 32:19]
  wire [63:0] idu_io_dataEx_dOut2; // @[riscv.scala 32:19]
  wire [63:0] idu_io_dataEx_dIn; // @[riscv.scala 32:19]
  wire [4:0] idu_io_rdOut; // @[riscv.scala 32:19]
  wire [4:0] idu_io_rdIn; // @[riscv.scala 32:19]
  wire [4:0] idu_io_rs1; // @[riscv.scala 32:19]
  wire [4:0] idu_io_rs2; // @[riscv.scala 32:19]
  wire [4:0] idu_io_rsWB; // @[riscv.scala 32:19]
  wire [63:0] idu_io_dOutWB; // @[riscv.scala 32:19]
  wire  idu_block1; // @[riscv.scala 32:19]
  wire  idu_block23; // @[riscv.scala 32:19]
  wire  exu_clock; // @[riscv.scala 33:19]
  wire  exu_reset; // @[riscv.scala 33:19]
  wire [1:0] exu_io_AluSrc1; // @[riscv.scala 33:19]
  wire [1:0] exu_io_AluSrc2; // @[riscv.scala 33:19]
  wire [4:0] exu_io_ALUCtrl; // @[riscv.scala 33:19]
  wire  exu_io_dnpcSrc; // @[riscv.scala 33:19]
  wire [1:0] exu_io_ResultSrc; // @[riscv.scala 33:19]
  wire [2:0] exu_io_memReadNum; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataId_imme; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataId_dOut1; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataId_dOut2; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataId_dIn; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataOut_ALUResOut; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataOut_wdata; // @[riscv.scala 33:19]
  wire [63:0] exu_io_dataOut_rdata; // @[riscv.scala 33:19]
  wire  exu_io_brTake; // @[riscv.scala 33:19]
  wire [31:0] exu_io_pc; // @[riscv.scala 33:19]
  wire [31:0] exu_io_snpc; // @[riscv.scala 33:19]
  wire [31:0] exu_io_dnpc; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrrwen; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrswen; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrrsien; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrrcien; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrrcen; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_csrrwien; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_ecall; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_rfen; // @[riscv.scala 33:19]
  wire  exu_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 33:19]
  wire [4:0] exu_io_uimm; // @[riscv.scala 33:19]
  wire [63:0] exu_io_aluResIn; // @[riscv.scala 33:19]
  wire [1:0] exu_io_forwardA; // @[riscv.scala 33:19]
  wire [1:0] exu_io_forwardB; // @[riscv.scala 33:19]
  wire [63:0] exu_io_aluRes1; // @[riscv.scala 33:19]
  wire [63:0] exu_io_aluRes3; // @[riscv.scala 33:19]
  wire  exu_intrTimeCnt_0; // @[riscv.scala 33:19]
  wire  exu_startTimeCnt; // @[riscv.scala 33:19]
  wire  exu_block1; // @[riscv.scala 33:19]
  wire  exu_block23; // @[riscv.scala 33:19]
  wire  hazardu_io_regEnEXMEM; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rdEXMEM; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rs1IDEX; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rs2IDEX; // @[riscv.scala 34:23]
  wire  hazardu_io_regEnMEMWB; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rdMEMWB; // @[riscv.scala 34:23]
  wire  hazardu_io_regEnWBEND; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rdWBEND; // @[riscv.scala 34:23]
  wire [1:0] hazardu_io_forwardA; // @[riscv.scala 34:23]
  wire [1:0] hazardu_io_forwardB; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rs1IFID; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rs2IFID; // @[riscv.scala 34:23]
  wire [4:0] hazardu_io_rdIDEX; // @[riscv.scala 34:23]
  wire [1:0] hazardu_io_resSrc; // @[riscv.scala 34:23]
  wire  hazardu_io_loadHazard; // @[riscv.scala 34:23]
  wire  preBranchIns_clock; // @[riscv.scala 35:28]
  wire  preBranchIns_reset; // @[riscv.scala 35:28]
  wire  preBranchIns_io_exjump; // @[riscv.scala 35:28]
  wire [31:0] preBranchIns_io_ifpc; // @[riscv.scala 35:28]
  wire [31:0] preBranchIns_io_expc; // @[riscv.scala 35:28]
  wire [31:0] preBranchIns_io_exdpc; // @[riscv.scala 35:28]
  wire [31:0] preBranchIns_io_ifdnpc; // @[riscv.scala 35:28]
  wire  preBranchIns_io_ifjump; // @[riscv.scala 35:28]
  wire  preBranchIns_block1_0; // @[riscv.scala 35:28]
  wire  preBranchIns_block23_0; // @[riscv.scala 35:28]
  wire [31:0] memVGenInst_io_inst; // @[riscv.scala 56:28]
  wire  memVGenInst_io_valid; // @[riscv.scala 56:28]
  wire [31:0] ctrl_io_inst; // @[riscv.scala 68:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc1; // @[riscv.scala 68:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc2; // @[riscv.scala 68:20]
  wire [4:0] ctrl_io_CtrlS_ALUCtrl; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_memWriteM; // @[riscv.scala 68:20]
  wire [7:0] ctrl_io_CtrlS_memWriteMask; // @[riscv.scala 68:20]
  wire [2:0] ctrl_io_CtrlS_memReadNum; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_dnpcSrc; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_jump; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_branch; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_regEn; // @[riscv.scala 68:20]
  wire [1:0] ctrl_io_CtrlS_ResultSrc; // @[riscv.scala 68:20]
  wire  ctrl_io_CtrlS_fencei; // @[riscv.scala 68:20]
  wire [31:0] csrCtrl_io_inst; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwen; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrswen; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrsien; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcien; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcen; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwien; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_ecall; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_rfen; // @[riscv.scala 69:23]
  wire  csrCtrl_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 69:23]
  wire  difftest_v; // @[riscv.scala 383:24]
  wire  intrins_intr; // @[riscv.scala 389:23]
  wire  Ebpro_block; // @[riscv.scala 395:21]
  wire [31:0] Ebpro_inst; // @[riscv.scala 395:21]
  wire  skipinst_v; // @[riscv.scala 399:24]
  wire  block1_0 = exu_block1;
  wire  _T = ~block1_0; // @[riscv.scala 49:32]
  wire  _T_2 = ~io_instIO_ready; // @[riscv.scala 53:23]
  wire  _T_3 = _T_2; // @[riscv.scala 53:20]
  wire  block2 = _T_2; // @[riscv.scala 52:20 riscv.scala 53:10]
  reg [247:0] pipEX2MEMReg; // @[Reg.scala 27:20]
  wire  pipEX2MEMWire_valid = pipEX2MEMReg[46]; // @[riscv.scala 253:44]
  wire  _T_159 = ~io_dataIO_ready; // @[riscv.scala 268:36]
  wire  _T_160 = pipEX2MEMWire_valid & _T_159; // @[riscv.scala 268:33]
  wire  block3 = _T_160; // @[riscv.scala 267:20 riscv.scala 268:10]
  wire  _T_161 = _T_3 | block3; // @[riscv.scala 273:21]
  wire  block23 = _T_161; // @[riscv.scala 272:23 riscv.scala 273:11]
  wire  pipBlock = block1_0 | block23; // @[riscv.scala 375:22]
  wire  _T_8 = ~pipBlock; // @[riscv.scala 95:30]
  reg [365:0] _T_59; // @[Reg.scala 27:20]
  wire  pipID2ExWire_branch = _T_59[47]; // @[riscv.scala 170:41]
  wire  _T_203 = pipID2ExWire_branch & exu_io_brTake; // @[riscv.scala 330:51]
  wire  pipID2ExWire_jump = _T_59[48]; // @[riscv.scala 170:41]
  wire  _T_204 = _T_203 | pipID2ExWire_jump; // @[riscv.scala 330:69]
  reg [8:0] _T_96; // @[Reg.scala 27:20]
  wire  pipCSRRegWire_mepc2pc = _T_96[0]; // @[riscv.scala 211:41]
  wire  _T_205 = _T_204 | pipCSRRegWire_mepc2pc; // @[riscv.scala 330:90]
  wire  pipCSRRegWire_ecall = _T_96[2]; // @[riscv.scala 211:41]
  wire  dnpcTakenWithoutPreB = _T_205 | pipCSRRegWire_ecall; // @[riscv.scala 330:115]
  wire  _T_206 = ~dnpcTakenWithoutPreB; // @[riscv.scala 331:15]
  wire  pipID2ExWire_ifjump = _T_59[32]; // @[riscv.scala 170:41]
  wire  jump1 = _T_206 & pipID2ExWire_ifjump; // @[riscv.scala 331:37]
  wire [31:0] pipID2ExWire_ifdnpc = _T_59[31:0]; // @[riscv.scala 170:41]
  wire  _T_207 = exu_io_dnpc != pipID2ExWire_ifdnpc; // @[riscv.scala 332:52]
  wire  _T_208 = ~pipID2ExWire_ifjump; // @[riscv.scala 332:79]
  wire  _T_209 = _T_207 | _T_208; // @[riscv.scala 332:76]
  wire  jump2 = dnpcTakenWithoutPreB & _T_209; // @[riscv.scala 332:36]
  wire  _T_210 = jump1 | jump2; // @[riscv.scala 333:25]
  wire [31:0] pipID2ExWire_pc = _T_59[140:109]; // @[riscv.scala 170:41]
  wire  _T_211 = pipID2ExWire_pc != 32'h0; // @[riscv.scala 333:69]
  wire  _T_212 = intrTimeCnt_0 & _T_211; // @[riscv.scala 333:50]
  wire  _T_213 = _T_210 | _T_212; // @[riscv.scala 333:34]
  wire  pipID2ExWire_fencei = _T_59[33]; // @[riscv.scala 170:41]
  wire  pipFlashWire = _T_213 | pipID2ExWire_fencei; // @[riscv.scala 333:78]
  wire  _T_9 = pipFlashWire & _T_8; // @[riscv.scala 95:27]
  wire  _T_11 = _T_9 | reset; // @[riscv.scala 95:40]
  wire  _T_12 = ifu_io_pc != 32'h0; // @[riscv.scala 97:16]
  wire [129:0] _T_17 = {_T_12,ifu_io_instOut,ifu_io_pc,ifu_io_snpc,preBranchIns_io_ifjump,preBranchIns_io_ifdnpc}; // @[Cat.scala 29:58]
  wire  _T_18 = pipBlock | hazardu_io_loadHazard; // @[riscv.scala 103:24]
  wire  _T_19 = ~_T_18; // @[riscv.scala 103:13]
  reg [129:0] _T_20; // @[Reg.scala 27:20]
  wire [31:0] pipIF2IDWire_ifdnpc = _T_20[31:0]; // @[riscv.scala 105:41]
  wire  pipIF2IDWire_ifjump = _T_20[32]; // @[riscv.scala 105:41]
  wire [31:0] pipIF2IDWire_snpc = _T_20[64:33]; // @[riscv.scala 105:41]
  wire [31:0] pipIF2IDWire_pc = _T_20[96:65]; // @[riscv.scala 105:41]
  wire [31:0] pipIF2IDWire_inst = _T_20[128:97]; // @[riscv.scala 105:41]
  wire  pipIF2IDWire_cmd = _T_20[129]; // @[riscv.scala 105:41]
  wire  _T_29 = pipFlashWire | hazardu_io_loadHazard; // @[riscv.scala 140:28]
  wire  _T_31 = _T_29 & _T_8; // @[riscv.scala 140:54]
  wire  _T_33 = _T_31 | reset; // @[riscv.scala 140:67]
  wire [45:0] _T_38 = {ctrl_io_CtrlS_ResultSrc,idu_io_rs1,idu_io_rs2,ctrl_io_CtrlS_fencei,pipIF2IDWire_ifjump,pipIF2IDWire_ifdnpc}; // @[Cat.scala 29:58]
  wire [58:0] _T_44 = {ctrl_io_CtrlS_memWriteMask,ctrl_io_CtrlS_memWriteM,ctrl_io_CtrlS_dnpcSrc,ctrl_io_CtrlS_jump,ctrl_io_CtrlS_branch,ctrl_io_CtrlS_regEn,_T_38}; // @[Cat.scala 29:58]
  wire [17:0] _T_49 = {idu_io_rdOut,ctrl_io_CtrlS_ALUCtrl,ctrl_io_CtrlS_AluSrc1,ctrl_io_CtrlS_AluSrc2,ctrl_io_CtrlS_memReadNum,memVGenInst_io_valid}; // @[Cat.scala 29:58]
  wire [365:0] _T_57 = {pipIF2IDWire_cmd,pipIF2IDWire_inst,idu_io_dataEx_imme,idu_io_dataEx_dOut1,idu_io_dataEx_dOut2,pipIF2IDWire_pc,pipIF2IDWire_snpc,_T_49,_T_44}; // @[Cat.scala 29:58]
  wire [1:0] pipID2ExWire_resultSrc = _T_59[45:44]; // @[riscv.scala 170:41]
  wire  pipID2ExWire_regEn = _T_59[46]; // @[riscv.scala 170:41]
  wire  pipID2ExWire_memWriteM = _T_59[50]; // @[riscv.scala 170:41]
  wire [7:0] pipID2ExWire_mask = _T_59[58:51]; // @[riscv.scala 170:41]
  wire  pipID2ExWire_valid = _T_59[59]; // @[riscv.scala 170:41]
  wire [2:0] pipID2ExWire_memReadNum = _T_59[62:60]; // @[riscv.scala 170:41]
  wire [4:0] pipID2ExWire_rd = _T_59[76:72]; // @[riscv.scala 170:41]
  wire [31:0] pipID2ExWire_snpc = _T_59[108:77]; // @[riscv.scala 170:41]
  wire [31:0] pipID2ExWire_inst = _T_59[364:333]; // @[riscv.scala 170:41]
  wire  pipID2ExWire_cmd = _T_59[365]; // @[riscv.scala 170:41]
  wire [8:0] _T_94 = {csrCtrl_io_CSRCtrlIf_csrrwen,csrCtrl_io_CSRCtrlIf_csrswen,csrCtrl_io_CSRCtrlIf_csrrsien,csrCtrl_io_CSRCtrlIf_csrrcien,csrCtrl_io_CSRCtrlIf_csrrcen,csrCtrl_io_CSRCtrlIf_csrrwien,csrCtrl_io_CSRCtrlIf_ecall,csrCtrl_io_CSRCtrlIf_rfen,csrCtrl_io_CSRCtrlIf_mepc2pc}; // @[Cat.scala 29:58]
  wire  pipCSRRegWire_rfen = _T_96[1]; // @[riscv.scala 211:41]
  wire  _T_110 = pipID2ExWire_regEn | pipCSRRegWire_rfen; // @[riscv.scala 247:21]
  wire [45:0] _T_118 = {pipID2ExWire_mask,pipID2ExWire_memWriteM,_T_110,pipID2ExWire_resultSrc,pipID2ExWire_pc,pipID2ExWire_fencei,_T_212}; // @[Cat.scala 29:58]
  wire [247:0] _T_126 = {pipID2ExWire_cmd,pipID2ExWire_inst,exu_io_dataOut_ALUResOut,exu_io_dataOut_wdata,pipID2ExWire_snpc,pipID2ExWire_rd,pipID2ExWire_memReadNum,pipID2ExWire_valid,_T_118}; // @[Cat.scala 29:58]
  wire  pipEX2MEMWire_intr = pipEX2MEMReg[0]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_fencei = pipEX2MEMReg[1]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_pc = pipEX2MEMReg[33:2]; // @[riscv.scala 253:44]
  wire [1:0] pipEX2MEMWire_ResultSrc = pipEX2MEMReg[35:34]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_regEn = pipEX2MEMReg[36]; // @[riscv.scala 253:44]
  wire [7:0] pipEX2MEMWire_mask = pipEX2MEMReg[45:38]; // @[riscv.scala 253:44]
  wire [2:0] pipEX2MEMWire_memReadNum = pipEX2MEMReg[49:47]; // @[riscv.scala 253:44]
  wire [4:0] pipEX2MEMWire_rd = pipEX2MEMReg[54:50]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_snpc = pipEX2MEMReg[86:55]; // @[riscv.scala 253:44]
  wire [63:0] pipEX2MEMWire_writeDataM = pipEX2MEMReg[150:87]; // @[riscv.scala 253:44]
  wire [63:0] pipEX2MEMWire_ALURes = pipEX2MEMReg[214:151]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_inst = pipEX2MEMReg[246:215]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_cmd = pipEX2MEMReg[247]; // @[riscv.scala 253:44]
  wire [14:0] _GEN_7 = {{7'd0}, pipEX2MEMWire_mask}; // @[riscv.scala 256:40]
  wire [14:0] _T_146 = _GEN_7 << pipEX2MEMWire_ALURes[2:0]; // @[riscv.scala 256:40]
  wire [3:0] _GEN_8 = {{1'd0}, pipEX2MEMWire_ALURes[2:0]}; // @[riscv.scala 261:78]
  wire [6:0] _T_149 = _GEN_8 * 4'h8; // @[riscv.scala 261:78]
  wire [190:0] _GEN_9 = {{127'd0}, pipEX2MEMWire_writeDataM}; // @[riscv.scala 261:50]
  wire [190:0] _T_150 = _GEN_9 << _T_149; // @[riscv.scala 261:50]
  wire  _T_153 = pipEX2MEMWire_ResultSrc == 2'h0; // @[riscv.scala 263:49]
  wire  _T_155 = pipEX2MEMWire_ALURes < 64'h80000000; // @[riscv.scala 265:59]
  wire  _T_156 = pipEX2MEMWire_ALURes > 64'h8fffffff; // @[riscv.scala 265:95]
  wire  _T_157 = _T_155 | _T_156; // @[riscv.scala 265:71]
  wire  _T_158 = pipEX2MEMWire_valid & _T_157; // @[riscv.scala 265:34]
  wire  skip = _T_158 | pipEX2MEMWire_fencei; // @[riscv.scala 265:109]
  wire  jud = pipEX2MEMWire_pc == 32'h0; // @[riscv.scala 278:29]
  reg [173:0] pipMEM2WBReg; // @[Reg.scala 27:20]
  wire [31:0] pipMEM2WBWire_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 293:44]
  wire [31:0] _T_186 = pipMEM2WBWire_pc + 32'h4; // @[riscv.scala 294:42]
  wire [31:0] npcsend = jud ? _T_186 : pipEX2MEMWire_pc; // @[riscv.scala 294:17]
  wire [36:0] _T_165 = {pipEX2MEMWire_regEn,pipEX2MEMWire_ResultSrc,npcsend,pipEX2MEMWire_intr,skip}; // @[Cat.scala 29:58]
  wire [173:0] _T_171 = {pipEX2MEMWire_cmd,pipEX2MEMWire_inst,pipEX2MEMWire_ALURes,pipEX2MEMWire_rd,pipEX2MEMWire_snpc,pipEX2MEMWire_memReadNum,_T_165}; // @[Cat.scala 29:58]
  wire  pipMEM2WBWire_intr = pipMEM2WBReg[1]; // @[riscv.scala 293:44]
  wire  pipMEM2WBWire_regEn = pipMEM2WBReg[36]; // @[riscv.scala 293:44]
  wire [4:0] pipMEM2WBWire_rd = pipMEM2WBReg[76:72]; // @[riscv.scala 293:44]
  wire [63:0] pipMEM2WBWire_ALURes = pipMEM2WBReg[140:77]; // @[riscv.scala 293:44]
  wire [31:0] pipMEM2WBWire_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 293:44]
  wire  pipMEM2WBWire_cmd = pipMEM2WBReg[173]; // @[riscv.scala 293:44]
  reg [63:0] _T_189; // @[Reg.scala 27:20]
  wire [3:0] _GEN_10 = {{1'd0}, pipMEM2WBWire_ALURes[2:0]}; // @[riscv.scala 302:100]
  wire [6:0] _T_191 = _GEN_10 * 4'h8; // @[riscv.scala 302:100]
  wire [69:0] _T_195 = {pipMEM2WBWire_rd,pipMEM2WBWire_regEn,pipMEM2WBWire_inst,pipMEM2WBWire_pc}; // @[Cat.scala 29:58]
  reg [69:0] _T_197; // @[Reg.scala 27:20]
  wire [31:0] _T_223 = jump2 ? exu_io_dnpc : preBranchIns_io_ifdnpc; // @[riscv.scala 345:12]
  wire [31:0] _T_224 = jump1 ? pipID2ExWire_snpc : _T_223; // @[riscv.scala 342:10]
  wire [31:0] _T_225 = pipID2ExWire_fencei ? pipID2ExWire_snpc : _T_224; // @[riscv.scala 339:8]
  wire  _T_228 = ~intrTimeCnt_0; // @[riscv.scala 378:36]
  wire  _T_229 = pipID2ExWire_fencei & _T_228; // @[riscv.scala 378:33]
  wire  _T_231 = _T_229 & _T_8; // @[riscv.scala 378:49]
  wire  hazardPCBlock = hazardu_io_loadHazard; // @[riscv.scala 371:27 riscv.scala 372:17]
  wire  fencei = _T_231; // @[riscv.scala 377:20 riscv.scala 378:10]
  iFetch ifu ( // @[riscv.scala 31:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_instIn(ifu_io_instIn),
    .io_instOut(ifu_io_instOut),
    .io_pc(ifu_io_pc),
    .io_snpc(ifu_io_snpc),
    .io_dnpc(ifu_io_dnpc),
    .io_jump(ifu_io_jump),
    .intrTimeCnt_0(ifu_intrTimeCnt_0),
    .hazardPCBlock_0(ifu_hazardPCBlock_0),
    .block1_0(ifu_block1_0),
    .block23_0(ifu_block23_0)
  );
  iDecode idu ( // @[riscv.scala 32:19]
    .clock(idu_clock),
    .io_pc(idu_io_pc),
    .io_inst(idu_io_inst),
    .io_regEn(idu_io_regEn),
    .io_dataEx_imme(idu_io_dataEx_imme),
    .io_dataEx_dOut1(idu_io_dataEx_dOut1),
    .io_dataEx_dOut2(idu_io_dataEx_dOut2),
    .io_dataEx_dIn(idu_io_dataEx_dIn),
    .io_rdOut(idu_io_rdOut),
    .io_rdIn(idu_io_rdIn),
    .io_rs1(idu_io_rs1),
    .io_rs2(idu_io_rs2),
    .io_rsWB(idu_io_rsWB),
    .io_dOutWB(idu_io_dOutWB),
    .block1(idu_block1),
    .block23(idu_block23)
  );
  execute exu ( // @[riscv.scala 33:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_AluSrc1(exu_io_AluSrc1),
    .io_AluSrc2(exu_io_AluSrc2),
    .io_ALUCtrl(exu_io_ALUCtrl),
    .io_dnpcSrc(exu_io_dnpcSrc),
    .io_ResultSrc(exu_io_ResultSrc),
    .io_memReadNum(exu_io_memReadNum),
    .io_dataId_imme(exu_io_dataId_imme),
    .io_dataId_dOut1(exu_io_dataId_dOut1),
    .io_dataId_dOut2(exu_io_dataId_dOut2),
    .io_dataId_dIn(exu_io_dataId_dIn),
    .io_dataOut_ALUResOut(exu_io_dataOut_ALUResOut),
    .io_dataOut_wdata(exu_io_dataOut_wdata),
    .io_dataOut_rdata(exu_io_dataOut_rdata),
    .io_brTake(exu_io_brTake),
    .io_pc(exu_io_pc),
    .io_snpc(exu_io_snpc),
    .io_dnpc(exu_io_dnpc),
    .io_CSRCtrlIf_csrrwen(exu_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(exu_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(exu_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(exu_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(exu_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(exu_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(exu_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(exu_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(exu_io_CSRCtrlIf_mepc2pc),
    .io_uimm(exu_io_uimm),
    .io_aluResIn(exu_io_aluResIn),
    .io_forwardA(exu_io_forwardA),
    .io_forwardB(exu_io_forwardB),
    .io_aluRes1(exu_io_aluRes1),
    .io_aluRes3(exu_io_aluRes3),
    .intrTimeCnt_0(exu_intrTimeCnt_0),
    .startTimeCnt(exu_startTimeCnt),
    .block1(exu_block1),
    .block23(exu_block23)
  );
  hazard hazardu ( // @[riscv.scala 34:23]
    .io_regEnEXMEM(hazardu_io_regEnEXMEM),
    .io_rdEXMEM(hazardu_io_rdEXMEM),
    .io_rs1IDEX(hazardu_io_rs1IDEX),
    .io_rs2IDEX(hazardu_io_rs2IDEX),
    .io_regEnMEMWB(hazardu_io_regEnMEMWB),
    .io_rdMEMWB(hazardu_io_rdMEMWB),
    .io_regEnWBEND(hazardu_io_regEnWBEND),
    .io_rdWBEND(hazardu_io_rdWBEND),
    .io_forwardA(hazardu_io_forwardA),
    .io_forwardB(hazardu_io_forwardB),
    .io_rs1IFID(hazardu_io_rs1IFID),
    .io_rs2IFID(hazardu_io_rs2IFID),
    .io_rdIDEX(hazardu_io_rdIDEX),
    .io_resSrc(hazardu_io_resSrc),
    .io_loadHazard(hazardu_io_loadHazard)
  );
  preBranch preBranchIns ( // @[riscv.scala 35:28]
    .clock(preBranchIns_clock),
    .reset(preBranchIns_reset),
    .io_exjump(preBranchIns_io_exjump),
    .io_ifpc(preBranchIns_io_ifpc),
    .io_expc(preBranchIns_io_expc),
    .io_exdpc(preBranchIns_io_exdpc),
    .io_ifdnpc(preBranchIns_io_ifdnpc),
    .io_ifjump(preBranchIns_io_ifjump),
    .block1_0(preBranchIns_block1_0),
    .block23_0(preBranchIns_block23_0)
  );
  memVGen memVGenInst ( // @[riscv.scala 56:28]
    .io_inst(memVGenInst_io_inst),
    .io_valid(memVGenInst_io_valid)
  );
  CtrlUnit ctrl ( // @[riscv.scala 68:20]
    .io_inst(ctrl_io_inst),
    .io_CtrlS_AluSrc1(ctrl_io_CtrlS_AluSrc1),
    .io_CtrlS_AluSrc2(ctrl_io_CtrlS_AluSrc2),
    .io_CtrlS_ALUCtrl(ctrl_io_CtrlS_ALUCtrl),
    .io_CtrlS_memWriteM(ctrl_io_CtrlS_memWriteM),
    .io_CtrlS_memWriteMask(ctrl_io_CtrlS_memWriteMask),
    .io_CtrlS_memReadNum(ctrl_io_CtrlS_memReadNum),
    .io_CtrlS_dnpcSrc(ctrl_io_CtrlS_dnpcSrc),
    .io_CtrlS_jump(ctrl_io_CtrlS_jump),
    .io_CtrlS_branch(ctrl_io_CtrlS_branch),
    .io_CtrlS_regEn(ctrl_io_CtrlS_regEn),
    .io_CtrlS_ResultSrc(ctrl_io_CtrlS_ResultSrc),
    .io_CtrlS_fencei(ctrl_io_CtrlS_fencei)
  );
  csrCtrl csrCtrl ( // @[riscv.scala 69:23]
    .io_inst(csrCtrl_io_inst),
    .io_CSRCtrlIf_csrrwen(csrCtrl_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(csrCtrl_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(csrCtrl_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(csrCtrl_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(csrCtrl_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(csrCtrl_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(csrCtrl_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(csrCtrl_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(csrCtrl_io_CSRCtrlIf_mepc2pc)
  );
  difftest difftest ( // @[riscv.scala 383:24]
    .v(difftest_v)
  );
  intr intrins ( // @[riscv.scala 389:23]
    .intr(intrins_intr)
  );
  ebProbe Ebpro ( // @[riscv.scala 395:21]
    .block(Ebpro_block),
    .inst(Ebpro_inst)
  );
  skip skipinst ( // @[riscv.scala 399:24]
    .v(skipinst_v)
  );
  assign io_instIO_valid = ~block1_0; // @[riscv.scala 49:19]
  assign io_instIO_addr = ifu_io_pc; // @[riscv.scala 88:18]
  assign io_dataIO_valid = pipEX2MEMWire_valid & _T; // @[riscv.scala 262:19]
  assign io_dataIO_data_write = _T_150[63:0]; // @[riscv.scala 261:23]
  assign io_dataIO_wen = pipEX2MEMReg[37]; // @[riscv.scala 257:17]
  assign io_dataIO_addr = pipEX2MEMWire_ALURes[31:0]; // @[riscv.scala 259:18]
  assign io_dataIO_rsize = pipEX2MEMWire_memReadNum[1:0]; // @[riscv.scala 260:19]
  assign io_dataIO_mask = _T_146[7:0]; // @[riscv.scala 256:18]
  assign startTimeCnt = exu_startTimeCnt;
  assign block2_0 = _T_3;
  assign fencei_0 = fencei;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_instIn = ifu_io_pc[2] ? io_instIO_data_read[63:32] : io_instIO_data_read[31:0]; // @[riscv.scala 87:17]
  assign ifu_io_dnpc = _T_212 ? exu_io_dnpc : _T_225; // @[riscv.scala 336:15]
  assign ifu_io_jump = pipFlashWire | preBranchIns_io_ifjump; // @[riscv.scala 335:15]
  assign ifu_intrTimeCnt_0 = intrTimeCnt_0;
  assign ifu_hazardPCBlock_0 = hazardPCBlock;
  assign ifu_block1_0 = exu_block1;
  assign ifu_block23_0 = block23;
  assign idu_clock = clock;
  assign idu_io_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 305:13]
  assign idu_io_inst = _T_20[128:97]; // @[riscv.scala 110:17]
  assign idu_io_regEn = pipMEM2WBReg[36]; // @[riscv.scala 299:16]
  assign idu_io_dataEx_dIn = exu_io_dataId_dIn; // @[riscv.scala 303:21]
  assign idu_io_rdIn = pipMEM2WBReg[76:72]; // @[riscv.scala 296:15]
  assign idu_io_rsWB = _T_197[69:65]; // @[riscv.scala 325:15]
  assign idu_block1 = exu_block1;
  assign idu_block23 = block23;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_AluSrc1 = _T_59[66:65]; // @[riscv.scala 179:20]
  assign exu_io_AluSrc2 = _T_59[64:63]; // @[riscv.scala 180:20]
  assign exu_io_ALUCtrl = _T_59[71:67]; // @[riscv.scala 178:19]
  assign exu_io_dnpcSrc = _T_59[49]; // @[riscv.scala 185:20]
  assign exu_io_ResultSrc = pipMEM2WBReg[35:34]; // @[riscv.scala 300:20]
  assign exu_io_memReadNum = pipMEM2WBReg[39:37]; // @[riscv.scala 298:21]
  assign exu_io_dataId_imme = _T_59[332:269]; // @[riscv.scala 172:24]
  assign exu_io_dataId_dOut1 = _T_59[268:205]; // @[riscv.scala 173:25]
  assign exu_io_dataId_dOut2 = _T_59[204:141]; // @[riscv.scala 174:25]
  assign exu_io_dataOut_rdata = _T_189 >> _T_191; // @[riscv.scala 302:24]
  assign exu_io_pc = _T_59[140:109]; // @[riscv.scala 175:15]
  assign exu_io_snpc = pipMEM2WBReg[71:40]; // @[riscv.scala 297:15]
  assign exu_io_CSRCtrlIf_csrrwen = _T_96[8]; // @[riscv.scala 212:30]
  assign exu_io_CSRCtrlIf_csrswen = _T_96[7]; // @[riscv.scala 213:30]
  assign exu_io_CSRCtrlIf_csrrsien = _T_96[6]; // @[riscv.scala 214:31]
  assign exu_io_CSRCtrlIf_csrrcien = _T_96[5]; // @[riscv.scala 215:31]
  assign exu_io_CSRCtrlIf_csrrcen = _T_96[4]; // @[riscv.scala 216:30]
  assign exu_io_CSRCtrlIf_csrrwien = _T_96[3]; // @[riscv.scala 217:31]
  assign exu_io_CSRCtrlIf_ecall = _T_96[2]; // @[riscv.scala 218:28]
  assign exu_io_CSRCtrlIf_rfen = _T_96[1]; // @[riscv.scala 219:27]
  assign exu_io_CSRCtrlIf_mepc2pc = _T_96[0]; // @[riscv.scala 221:30]
  assign exu_io_uimm = _T_59[43:39]; // @[riscv.scala 222:17]
  assign exu_io_aluResIn = pipMEM2WBReg[140:77]; // @[riscv.scala 295:19]
  assign exu_io_forwardA = hazardu_io_forwardA; // @[riscv.scala 362:19]
  assign exu_io_forwardB = hazardu_io_forwardB; // @[riscv.scala 363:19]
  assign exu_io_aluRes1 = _T_153 ? pipEX2MEMWire_ALURes : {{32'd0}, pipEX2MEMWire_snpc}; // @[riscv.scala 263:18]
  assign exu_io_aluRes3 = idu_io_dOutWB; // @[riscv.scala 326:18]
  assign exu_intrTimeCnt_0 = intrTimeCnt_0;
  assign exu_block23 = block23;
  assign hazardu_io_regEnEXMEM = pipEX2MEMReg[36]; // @[riscv.scala 355:25]
  assign hazardu_io_rdEXMEM = pipEX2MEMReg[54:50]; // @[riscv.scala 356:22]
  assign hazardu_io_rs1IDEX = _T_59[43:39]; // @[riscv.scala 192:24]
  assign hazardu_io_rs2IDEX = _T_59[38:34]; // @[riscv.scala 193:24]
  assign hazardu_io_regEnMEMWB = pipMEM2WBReg[36]; // @[riscv.scala 357:25]
  assign hazardu_io_rdMEMWB = pipMEM2WBReg[76:72]; // @[riscv.scala 358:22]
  assign hazardu_io_regEnWBEND = _T_197[64]; // @[riscv.scala 359:25]
  assign hazardu_io_rdWBEND = _T_197[69:65]; // @[riscv.scala 360:22]
  assign hazardu_io_rs1IFID = idu_io_rs1; // @[riscv.scala 366:22]
  assign hazardu_io_rs2IFID = idu_io_rs2; // @[riscv.scala 367:22]
  assign hazardu_io_rdIDEX = _T_59[76:72]; // @[riscv.scala 368:21]
  assign hazardu_io_resSrc = _T_59[45:44]; // @[riscv.scala 369:21]
  assign preBranchIns_clock = clock;
  assign preBranchIns_reset = reset;
  assign preBranchIns_io_exjump = _T_205 | pipCSRRegWire_ecall; // @[riscv.scala 548:26]
  assign preBranchIns_io_ifpc = ifu_io_pc; // @[riscv.scala 547:24]
  assign preBranchIns_io_expc = _T_59[140:109]; // @[riscv.scala 549:24]
  assign preBranchIns_io_exdpc = exu_io_dnpc; // @[riscv.scala 550:25]
  assign preBranchIns_block1_0 = exu_block1;
  assign preBranchIns_block23_0 = block23;
  assign memVGenInst_io_inst = _T_20[128:97]; // @[riscv.scala 107:25]
  assign ctrl_io_inst = _T_20[128:97]; // @[riscv.scala 109:18]
  assign csrCtrl_io_inst = _T_20[128:97]; // @[riscv.scala 108:21]
  assign difftest_v = pipMEM2WBWire_cmd & _T_8; // @[riscv.scala 384:17]
  assign intrins_intr = pipMEM2WBWire_intr & _T_8; // @[riscv.scala 390:19]
  assign Ebpro_block = block1_0 | block23; // @[riscv.scala 397:18]
  assign Ebpro_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 396:17]
  assign skipinst_v = pipMEM2WBReg[0]; // @[riscv.scala 400:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  pipEX2MEMReg = _RAND_0[247:0];
  _RAND_1 = {12{`RANDOM}};
  _T_59 = _RAND_1[365:0];
  _RAND_2 = {1{`RANDOM}};
  _T_96 = _RAND_2[8:0];
  _RAND_3 = {5{`RANDOM}};
  _T_20 = _RAND_3[129:0];
  _RAND_4 = {6{`RANDOM}};
  pipMEM2WBReg = _RAND_4[173:0];
  _RAND_5 = {2{`RANDOM}};
  _T_189 = _RAND_5[63:0];
  _RAND_6 = {3{`RANDOM}};
  _T_197 = _RAND_6[69:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pipEX2MEMReg <= 248'h0;
    end else if (_T_8) begin
      if (_T_212) begin
        pipEX2MEMReg <= 248'h1;
      end else begin
        pipEX2MEMReg <= _T_126;
      end
    end
    if (_T_33) begin
      _T_59 <= 366'h0;
    end else if (_T_8) begin
      _T_59 <= _T_57;
    end
    if (_T_33) begin
      _T_96 <= 9'h0;
    end else if (_T_8) begin
      _T_96 <= _T_94;
    end
    if (_T_11) begin
      _T_20 <= 130'h0;
    end else if (_T_19) begin
      _T_20 <= _T_17;
    end
    if (reset) begin
      pipMEM2WBReg <= 174'h0;
    end else if (_T_8) begin
      pipMEM2WBReg <= _T_171;
    end
    if (reset) begin
      _T_189 <= 64'h0;
    end else if (_T_8) begin
      _T_189 <= io_dataIO_data_read;
    end
    if (reset) begin
      _T_197 <= 70'h0;
    end else if (_T_8) begin
      _T_197 <= _T_195;
    end
  end
endmodule
module Icache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output [31:0]  io_cacheOut_w_addr_o,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [31:0]  io_cacheIn_addr,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          updataICache_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] offset = io_cacheIn_addr[3:0]; // @[Cache.scala 27:31]
  wire [5:0] index = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  wire [21:0] tag = io_cacheIn_addr[31:10]; // @[Cache.scala 29:28]
  reg  cacheState; // @[Cache.scala 32:27]
  wire  _T_253 = 6'h3f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_63_0; // @[Reg.scala 27:20]
  wire  _T_251 = 6'h3e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_62_0; // @[Reg.scala 27:20]
  wire  _T_249 = 6'h3d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_61_0; // @[Reg.scala 27:20]
  wire  _T_247 = 6'h3c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_60_0; // @[Reg.scala 27:20]
  wire  _T_245 = 6'h3b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_59_0; // @[Reg.scala 27:20]
  wire  _T_243 = 6'h3a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_58_0; // @[Reg.scala 27:20]
  wire  _T_241 = 6'h39 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_57_0; // @[Reg.scala 27:20]
  wire  _T_239 = 6'h38 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_56_0; // @[Reg.scala 27:20]
  wire  _T_237 = 6'h37 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_55_0; // @[Reg.scala 27:20]
  wire  _T_235 = 6'h36 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_54_0; // @[Reg.scala 27:20]
  wire  _T_233 = 6'h35 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_53_0; // @[Reg.scala 27:20]
  wire  _T_231 = 6'h34 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_52_0; // @[Reg.scala 27:20]
  wire  _T_229 = 6'h33 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_51_0; // @[Reg.scala 27:20]
  wire  _T_227 = 6'h32 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_50_0; // @[Reg.scala 27:20]
  wire  _T_225 = 6'h31 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_49_0; // @[Reg.scala 27:20]
  wire  _T_223 = 6'h30 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_48_0; // @[Reg.scala 27:20]
  wire  _T_221 = 6'h2f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_47_0; // @[Reg.scala 27:20]
  wire  _T_219 = 6'h2e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_46_0; // @[Reg.scala 27:20]
  wire  _T_217 = 6'h2d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_45_0; // @[Reg.scala 27:20]
  wire  _T_215 = 6'h2c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_44_0; // @[Reg.scala 27:20]
  wire  _T_213 = 6'h2b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_43_0; // @[Reg.scala 27:20]
  wire  _T_211 = 6'h2a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_42_0; // @[Reg.scala 27:20]
  wire  _T_209 = 6'h29 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_41_0; // @[Reg.scala 27:20]
  wire  _T_207 = 6'h28 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_40_0; // @[Reg.scala 27:20]
  wire  _T_205 = 6'h27 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_39_0; // @[Reg.scala 27:20]
  wire  _T_203 = 6'h26 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_38_0; // @[Reg.scala 27:20]
  wire  _T_201 = 6'h25 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_37_0; // @[Reg.scala 27:20]
  wire  _T_199 = 6'h24 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_36_0; // @[Reg.scala 27:20]
  wire  _T_197 = 6'h23 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_35_0; // @[Reg.scala 27:20]
  wire  _T_195 = 6'h22 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_34_0; // @[Reg.scala 27:20]
  wire  _T_193 = 6'h21 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_33_0; // @[Reg.scala 27:20]
  wire  _T_191 = 6'h20 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_32_0; // @[Reg.scala 27:20]
  wire  _T_189 = 6'h1f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_31_0; // @[Reg.scala 27:20]
  wire  _T_187 = 6'h1e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_30_0; // @[Reg.scala 27:20]
  wire  _T_185 = 6'h1d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_29_0; // @[Reg.scala 27:20]
  wire  _T_183 = 6'h1c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_28_0; // @[Reg.scala 27:20]
  wire  _T_181 = 6'h1b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_27_0; // @[Reg.scala 27:20]
  wire  _T_179 = 6'h1a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_26_0; // @[Reg.scala 27:20]
  wire  _T_177 = 6'h19 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_25_0; // @[Reg.scala 27:20]
  wire  _T_175 = 6'h18 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_24_0; // @[Reg.scala 27:20]
  wire  _T_173 = 6'h17 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_23_0; // @[Reg.scala 27:20]
  wire  _T_171 = 6'h16 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_22_0; // @[Reg.scala 27:20]
  wire  _T_169 = 6'h15 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_21_0; // @[Reg.scala 27:20]
  wire  _T_167 = 6'h14 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_20_0; // @[Reg.scala 27:20]
  wire  _T_165 = 6'h13 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_19_0; // @[Reg.scala 27:20]
  wire  _T_163 = 6'h12 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_18_0; // @[Reg.scala 27:20]
  wire  _T_161 = 6'h11 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_17_0; // @[Reg.scala 27:20]
  wire  _T_159 = 6'h10 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_16_0; // @[Reg.scala 27:20]
  wire  _T_157 = 6'hf == index; // @[Mux.scala 80:60]
  reg  vArrayWire_15_0; // @[Reg.scala 27:20]
  wire  _T_155 = 6'he == index; // @[Mux.scala 80:60]
  reg  vArrayWire_14_0; // @[Reg.scala 27:20]
  wire  _T_153 = 6'hd == index; // @[Mux.scala 80:60]
  reg  vArrayWire_13_0; // @[Reg.scala 27:20]
  wire  _T_151 = 6'hc == index; // @[Mux.scala 80:60]
  reg  vArrayWire_12_0; // @[Reg.scala 27:20]
  wire  _T_149 = 6'hb == index; // @[Mux.scala 80:60]
  reg  vArrayWire_11_0; // @[Reg.scala 27:20]
  wire  _T_147 = 6'ha == index; // @[Mux.scala 80:60]
  reg  vArrayWire_10_0; // @[Reg.scala 27:20]
  wire  _T_145 = 6'h9 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_9_0; // @[Reg.scala 27:20]
  wire  _T_143 = 6'h8 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_8_0; // @[Reg.scala 27:20]
  wire  _T_141 = 6'h7 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_7_0; // @[Reg.scala 27:20]
  wire  _T_139 = 6'h6 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_6_0; // @[Reg.scala 27:20]
  wire  _T_137 = 6'h5 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_5_0; // @[Reg.scala 27:20]
  wire  _T_135 = 6'h4 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_4_0; // @[Reg.scala 27:20]
  wire  _T_133 = 6'h3 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_3_0; // @[Reg.scala 27:20]
  wire  _T_131 = 6'h2 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_2_0; // @[Reg.scala 27:20]
  wire  _T_129 = 6'h1 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_1_0; // @[Reg.scala 27:20]
  reg  vArrayWire_0_0; // @[Reg.scala 27:20]
  wire  _T_130_0 = _T_129 ? vArrayWire_1_0 : vArrayWire_0_0; // @[Mux.scala 80:57]
  wire  _T_132_0 = _T_131 ? vArrayWire_2_0 : _T_130_0; // @[Mux.scala 80:57]
  wire  _T_134_0 = _T_133 ? vArrayWire_3_0 : _T_132_0; // @[Mux.scala 80:57]
  wire  _T_136_0 = _T_135 ? vArrayWire_4_0 : _T_134_0; // @[Mux.scala 80:57]
  wire  _T_138_0 = _T_137 ? vArrayWire_5_0 : _T_136_0; // @[Mux.scala 80:57]
  wire  _T_140_0 = _T_139 ? vArrayWire_6_0 : _T_138_0; // @[Mux.scala 80:57]
  wire  _T_142_0 = _T_141 ? vArrayWire_7_0 : _T_140_0; // @[Mux.scala 80:57]
  wire  _T_144_0 = _T_143 ? vArrayWire_8_0 : _T_142_0; // @[Mux.scala 80:57]
  wire  _T_146_0 = _T_145 ? vArrayWire_9_0 : _T_144_0; // @[Mux.scala 80:57]
  wire  _T_148_0 = _T_147 ? vArrayWire_10_0 : _T_146_0; // @[Mux.scala 80:57]
  wire  _T_150_0 = _T_149 ? vArrayWire_11_0 : _T_148_0; // @[Mux.scala 80:57]
  wire  _T_152_0 = _T_151 ? vArrayWire_12_0 : _T_150_0; // @[Mux.scala 80:57]
  wire  _T_154_0 = _T_153 ? vArrayWire_13_0 : _T_152_0; // @[Mux.scala 80:57]
  wire  _T_156_0 = _T_155 ? vArrayWire_14_0 : _T_154_0; // @[Mux.scala 80:57]
  wire  _T_158_0 = _T_157 ? vArrayWire_15_0 : _T_156_0; // @[Mux.scala 80:57]
  wire  _T_160_0 = _T_159 ? vArrayWire_16_0 : _T_158_0; // @[Mux.scala 80:57]
  wire  _T_162_0 = _T_161 ? vArrayWire_17_0 : _T_160_0; // @[Mux.scala 80:57]
  wire  _T_164_0 = _T_163 ? vArrayWire_18_0 : _T_162_0; // @[Mux.scala 80:57]
  wire  _T_166_0 = _T_165 ? vArrayWire_19_0 : _T_164_0; // @[Mux.scala 80:57]
  wire  _T_168_0 = _T_167 ? vArrayWire_20_0 : _T_166_0; // @[Mux.scala 80:57]
  wire  _T_170_0 = _T_169 ? vArrayWire_21_0 : _T_168_0; // @[Mux.scala 80:57]
  wire  _T_172_0 = _T_171 ? vArrayWire_22_0 : _T_170_0; // @[Mux.scala 80:57]
  wire  _T_174_0 = _T_173 ? vArrayWire_23_0 : _T_172_0; // @[Mux.scala 80:57]
  wire  _T_176_0 = _T_175 ? vArrayWire_24_0 : _T_174_0; // @[Mux.scala 80:57]
  wire  _T_178_0 = _T_177 ? vArrayWire_25_0 : _T_176_0; // @[Mux.scala 80:57]
  wire  _T_180_0 = _T_179 ? vArrayWire_26_0 : _T_178_0; // @[Mux.scala 80:57]
  wire  _T_182_0 = _T_181 ? vArrayWire_27_0 : _T_180_0; // @[Mux.scala 80:57]
  wire  _T_184_0 = _T_183 ? vArrayWire_28_0 : _T_182_0; // @[Mux.scala 80:57]
  wire  _T_186_0 = _T_185 ? vArrayWire_29_0 : _T_184_0; // @[Mux.scala 80:57]
  wire  _T_188_0 = _T_187 ? vArrayWire_30_0 : _T_186_0; // @[Mux.scala 80:57]
  wire  _T_190_0 = _T_189 ? vArrayWire_31_0 : _T_188_0; // @[Mux.scala 80:57]
  wire  _T_192_0 = _T_191 ? vArrayWire_32_0 : _T_190_0; // @[Mux.scala 80:57]
  wire  _T_194_0 = _T_193 ? vArrayWire_33_0 : _T_192_0; // @[Mux.scala 80:57]
  wire  _T_196_0 = _T_195 ? vArrayWire_34_0 : _T_194_0; // @[Mux.scala 80:57]
  wire  _T_198_0 = _T_197 ? vArrayWire_35_0 : _T_196_0; // @[Mux.scala 80:57]
  wire  _T_200_0 = _T_199 ? vArrayWire_36_0 : _T_198_0; // @[Mux.scala 80:57]
  wire  _T_202_0 = _T_201 ? vArrayWire_37_0 : _T_200_0; // @[Mux.scala 80:57]
  wire  _T_204_0 = _T_203 ? vArrayWire_38_0 : _T_202_0; // @[Mux.scala 80:57]
  wire  _T_206_0 = _T_205 ? vArrayWire_39_0 : _T_204_0; // @[Mux.scala 80:57]
  wire  _T_208_0 = _T_207 ? vArrayWire_40_0 : _T_206_0; // @[Mux.scala 80:57]
  wire  _T_210_0 = _T_209 ? vArrayWire_41_0 : _T_208_0; // @[Mux.scala 80:57]
  wire  _T_212_0 = _T_211 ? vArrayWire_42_0 : _T_210_0; // @[Mux.scala 80:57]
  wire  _T_214_0 = _T_213 ? vArrayWire_43_0 : _T_212_0; // @[Mux.scala 80:57]
  wire  _T_216_0 = _T_215 ? vArrayWire_44_0 : _T_214_0; // @[Mux.scala 80:57]
  wire  _T_218_0 = _T_217 ? vArrayWire_45_0 : _T_216_0; // @[Mux.scala 80:57]
  wire  _T_220_0 = _T_219 ? vArrayWire_46_0 : _T_218_0; // @[Mux.scala 80:57]
  wire  _T_222_0 = _T_221 ? vArrayWire_47_0 : _T_220_0; // @[Mux.scala 80:57]
  wire  _T_224_0 = _T_223 ? vArrayWire_48_0 : _T_222_0; // @[Mux.scala 80:57]
  wire  _T_226_0 = _T_225 ? vArrayWire_49_0 : _T_224_0; // @[Mux.scala 80:57]
  wire  _T_228_0 = _T_227 ? vArrayWire_50_0 : _T_226_0; // @[Mux.scala 80:57]
  wire  _T_230_0 = _T_229 ? vArrayWire_51_0 : _T_228_0; // @[Mux.scala 80:57]
  wire  _T_232_0 = _T_231 ? vArrayWire_52_0 : _T_230_0; // @[Mux.scala 80:57]
  wire  _T_234_0 = _T_233 ? vArrayWire_53_0 : _T_232_0; // @[Mux.scala 80:57]
  wire  _T_236_0 = _T_235 ? vArrayWire_54_0 : _T_234_0; // @[Mux.scala 80:57]
  wire  _T_238_0 = _T_237 ? vArrayWire_55_0 : _T_236_0; // @[Mux.scala 80:57]
  wire  _T_240_0 = _T_239 ? vArrayWire_56_0 : _T_238_0; // @[Mux.scala 80:57]
  wire  _T_242_0 = _T_241 ? vArrayWire_57_0 : _T_240_0; // @[Mux.scala 80:57]
  wire  _T_244_0 = _T_243 ? vArrayWire_58_0 : _T_242_0; // @[Mux.scala 80:57]
  wire  _T_246_0 = _T_245 ? vArrayWire_59_0 : _T_244_0; // @[Mux.scala 80:57]
  wire  _T_248_0 = _T_247 ? vArrayWire_60_0 : _T_246_0; // @[Mux.scala 80:57]
  wire  _T_250_0 = _T_249 ? vArrayWire_61_0 : _T_248_0; // @[Mux.scala 80:57]
  wire  _T_252_0 = _T_251 ? vArrayWire_62_0 : _T_250_0; // @[Mux.scala 80:57]
  wire  vMuxOut_0 = _T_253 ? vArrayWire_63_0 : _T_252_0; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_0; // @[Reg.scala 27:20]
  wire [21:0] _T_5_0 = _T_129 ? tagArrayWire_1_0 : tagArrayWire_0_0; // @[Mux.scala 80:57]
  wire [21:0] _T_7_0 = _T_131 ? tagArrayWire_2_0 : _T_5_0; // @[Mux.scala 80:57]
  wire [21:0] _T_9_0 = _T_133 ? tagArrayWire_3_0 : _T_7_0; // @[Mux.scala 80:57]
  wire [21:0] _T_11_0 = _T_135 ? tagArrayWire_4_0 : _T_9_0; // @[Mux.scala 80:57]
  wire [21:0] _T_13_0 = _T_137 ? tagArrayWire_5_0 : _T_11_0; // @[Mux.scala 80:57]
  wire [21:0] _T_15_0 = _T_139 ? tagArrayWire_6_0 : _T_13_0; // @[Mux.scala 80:57]
  wire [21:0] _T_17_0 = _T_141 ? tagArrayWire_7_0 : _T_15_0; // @[Mux.scala 80:57]
  wire [21:0] _T_19_0 = _T_143 ? tagArrayWire_8_0 : _T_17_0; // @[Mux.scala 80:57]
  wire [21:0] _T_21_0 = _T_145 ? tagArrayWire_9_0 : _T_19_0; // @[Mux.scala 80:57]
  wire [21:0] _T_23_0 = _T_147 ? tagArrayWire_10_0 : _T_21_0; // @[Mux.scala 80:57]
  wire [21:0] _T_25_0 = _T_149 ? tagArrayWire_11_0 : _T_23_0; // @[Mux.scala 80:57]
  wire [21:0] _T_27_0 = _T_151 ? tagArrayWire_12_0 : _T_25_0; // @[Mux.scala 80:57]
  wire [21:0] _T_29_0 = _T_153 ? tagArrayWire_13_0 : _T_27_0; // @[Mux.scala 80:57]
  wire [21:0] _T_31_0 = _T_155 ? tagArrayWire_14_0 : _T_29_0; // @[Mux.scala 80:57]
  wire [21:0] _T_33_0 = _T_157 ? tagArrayWire_15_0 : _T_31_0; // @[Mux.scala 80:57]
  wire [21:0] _T_35_0 = _T_159 ? tagArrayWire_16_0 : _T_33_0; // @[Mux.scala 80:57]
  wire [21:0] _T_37_0 = _T_161 ? tagArrayWire_17_0 : _T_35_0; // @[Mux.scala 80:57]
  wire [21:0] _T_39_0 = _T_163 ? tagArrayWire_18_0 : _T_37_0; // @[Mux.scala 80:57]
  wire [21:0] _T_41_0 = _T_165 ? tagArrayWire_19_0 : _T_39_0; // @[Mux.scala 80:57]
  wire [21:0] _T_43_0 = _T_167 ? tagArrayWire_20_0 : _T_41_0; // @[Mux.scala 80:57]
  wire [21:0] _T_45_0 = _T_169 ? tagArrayWire_21_0 : _T_43_0; // @[Mux.scala 80:57]
  wire [21:0] _T_47_0 = _T_171 ? tagArrayWire_22_0 : _T_45_0; // @[Mux.scala 80:57]
  wire [21:0] _T_49_0 = _T_173 ? tagArrayWire_23_0 : _T_47_0; // @[Mux.scala 80:57]
  wire [21:0] _T_51_0 = _T_175 ? tagArrayWire_24_0 : _T_49_0; // @[Mux.scala 80:57]
  wire [21:0] _T_53_0 = _T_177 ? tagArrayWire_25_0 : _T_51_0; // @[Mux.scala 80:57]
  wire [21:0] _T_55_0 = _T_179 ? tagArrayWire_26_0 : _T_53_0; // @[Mux.scala 80:57]
  wire [21:0] _T_57_0 = _T_181 ? tagArrayWire_27_0 : _T_55_0; // @[Mux.scala 80:57]
  wire [21:0] _T_59_0 = _T_183 ? tagArrayWire_28_0 : _T_57_0; // @[Mux.scala 80:57]
  wire [21:0] _T_61_0 = _T_185 ? tagArrayWire_29_0 : _T_59_0; // @[Mux.scala 80:57]
  wire [21:0] _T_63_0 = _T_187 ? tagArrayWire_30_0 : _T_61_0; // @[Mux.scala 80:57]
  wire [21:0] _T_65_0 = _T_189 ? tagArrayWire_31_0 : _T_63_0; // @[Mux.scala 80:57]
  wire [21:0] _T_67_0 = _T_191 ? tagArrayWire_32_0 : _T_65_0; // @[Mux.scala 80:57]
  wire [21:0] _T_69_0 = _T_193 ? tagArrayWire_33_0 : _T_67_0; // @[Mux.scala 80:57]
  wire [21:0] _T_71_0 = _T_195 ? tagArrayWire_34_0 : _T_69_0; // @[Mux.scala 80:57]
  wire [21:0] _T_73_0 = _T_197 ? tagArrayWire_35_0 : _T_71_0; // @[Mux.scala 80:57]
  wire [21:0] _T_75_0 = _T_199 ? tagArrayWire_36_0 : _T_73_0; // @[Mux.scala 80:57]
  wire [21:0] _T_77_0 = _T_201 ? tagArrayWire_37_0 : _T_75_0; // @[Mux.scala 80:57]
  wire [21:0] _T_79_0 = _T_203 ? tagArrayWire_38_0 : _T_77_0; // @[Mux.scala 80:57]
  wire [21:0] _T_81_0 = _T_205 ? tagArrayWire_39_0 : _T_79_0; // @[Mux.scala 80:57]
  wire [21:0] _T_83_0 = _T_207 ? tagArrayWire_40_0 : _T_81_0; // @[Mux.scala 80:57]
  wire [21:0] _T_85_0 = _T_209 ? tagArrayWire_41_0 : _T_83_0; // @[Mux.scala 80:57]
  wire [21:0] _T_87_0 = _T_211 ? tagArrayWire_42_0 : _T_85_0; // @[Mux.scala 80:57]
  wire [21:0] _T_89_0 = _T_213 ? tagArrayWire_43_0 : _T_87_0; // @[Mux.scala 80:57]
  wire [21:0] _T_91_0 = _T_215 ? tagArrayWire_44_0 : _T_89_0; // @[Mux.scala 80:57]
  wire [21:0] _T_93_0 = _T_217 ? tagArrayWire_45_0 : _T_91_0; // @[Mux.scala 80:57]
  wire [21:0] _T_95_0 = _T_219 ? tagArrayWire_46_0 : _T_93_0; // @[Mux.scala 80:57]
  wire [21:0] _T_97_0 = _T_221 ? tagArrayWire_47_0 : _T_95_0; // @[Mux.scala 80:57]
  wire [21:0] _T_99_0 = _T_223 ? tagArrayWire_48_0 : _T_97_0; // @[Mux.scala 80:57]
  wire [21:0] _T_101_0 = _T_225 ? tagArrayWire_49_0 : _T_99_0; // @[Mux.scala 80:57]
  wire [21:0] _T_103_0 = _T_227 ? tagArrayWire_50_0 : _T_101_0; // @[Mux.scala 80:57]
  wire [21:0] _T_105_0 = _T_229 ? tagArrayWire_51_0 : _T_103_0; // @[Mux.scala 80:57]
  wire [21:0] _T_107_0 = _T_231 ? tagArrayWire_52_0 : _T_105_0; // @[Mux.scala 80:57]
  wire [21:0] _T_109_0 = _T_233 ? tagArrayWire_53_0 : _T_107_0; // @[Mux.scala 80:57]
  wire [21:0] _T_111_0 = _T_235 ? tagArrayWire_54_0 : _T_109_0; // @[Mux.scala 80:57]
  wire [21:0] _T_113_0 = _T_237 ? tagArrayWire_55_0 : _T_111_0; // @[Mux.scala 80:57]
  wire [21:0] _T_115_0 = _T_239 ? tagArrayWire_56_0 : _T_113_0; // @[Mux.scala 80:57]
  wire [21:0] _T_117_0 = _T_241 ? tagArrayWire_57_0 : _T_115_0; // @[Mux.scala 80:57]
  wire [21:0] _T_119_0 = _T_243 ? tagArrayWire_58_0 : _T_117_0; // @[Mux.scala 80:57]
  wire [21:0] _T_121_0 = _T_245 ? tagArrayWire_59_0 : _T_119_0; // @[Mux.scala 80:57]
  wire [21:0] _T_123_0 = _T_247 ? tagArrayWire_60_0 : _T_121_0; // @[Mux.scala 80:57]
  wire [21:0] _T_125_0 = _T_249 ? tagArrayWire_61_0 : _T_123_0; // @[Mux.scala 80:57]
  wire [21:0] _T_127_0 = _T_251 ? tagArrayWire_62_0 : _T_125_0; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_0 = _T_253 ? tagArrayWire_63_0 : _T_127_0; // @[Mux.scala 80:57]
  wire  _T_254 = tagMuxOut_0 == tag; // @[Cache.scala 72:76]
  wire  hitArray_0 = vMuxOut_0 & _T_254; // @[Cache.scala 72:60]
  reg  vArrayWire_63_1; // @[Reg.scala 27:20]
  reg  vArrayWire_62_1; // @[Reg.scala 27:20]
  reg  vArrayWire_61_1; // @[Reg.scala 27:20]
  reg  vArrayWire_60_1; // @[Reg.scala 27:20]
  reg  vArrayWire_59_1; // @[Reg.scala 27:20]
  reg  vArrayWire_58_1; // @[Reg.scala 27:20]
  reg  vArrayWire_57_1; // @[Reg.scala 27:20]
  reg  vArrayWire_56_1; // @[Reg.scala 27:20]
  reg  vArrayWire_55_1; // @[Reg.scala 27:20]
  reg  vArrayWire_54_1; // @[Reg.scala 27:20]
  reg  vArrayWire_53_1; // @[Reg.scala 27:20]
  reg  vArrayWire_52_1; // @[Reg.scala 27:20]
  reg  vArrayWire_51_1; // @[Reg.scala 27:20]
  reg  vArrayWire_50_1; // @[Reg.scala 27:20]
  reg  vArrayWire_49_1; // @[Reg.scala 27:20]
  reg  vArrayWire_48_1; // @[Reg.scala 27:20]
  reg  vArrayWire_47_1; // @[Reg.scala 27:20]
  reg  vArrayWire_46_1; // @[Reg.scala 27:20]
  reg  vArrayWire_45_1; // @[Reg.scala 27:20]
  reg  vArrayWire_44_1; // @[Reg.scala 27:20]
  reg  vArrayWire_43_1; // @[Reg.scala 27:20]
  reg  vArrayWire_42_1; // @[Reg.scala 27:20]
  reg  vArrayWire_41_1; // @[Reg.scala 27:20]
  reg  vArrayWire_40_1; // @[Reg.scala 27:20]
  reg  vArrayWire_39_1; // @[Reg.scala 27:20]
  reg  vArrayWire_38_1; // @[Reg.scala 27:20]
  reg  vArrayWire_37_1; // @[Reg.scala 27:20]
  reg  vArrayWire_36_1; // @[Reg.scala 27:20]
  reg  vArrayWire_35_1; // @[Reg.scala 27:20]
  reg  vArrayWire_34_1; // @[Reg.scala 27:20]
  reg  vArrayWire_33_1; // @[Reg.scala 27:20]
  reg  vArrayWire_32_1; // @[Reg.scala 27:20]
  reg  vArrayWire_31_1; // @[Reg.scala 27:20]
  reg  vArrayWire_30_1; // @[Reg.scala 27:20]
  reg  vArrayWire_29_1; // @[Reg.scala 27:20]
  reg  vArrayWire_28_1; // @[Reg.scala 27:20]
  reg  vArrayWire_27_1; // @[Reg.scala 27:20]
  reg  vArrayWire_26_1; // @[Reg.scala 27:20]
  reg  vArrayWire_25_1; // @[Reg.scala 27:20]
  reg  vArrayWire_24_1; // @[Reg.scala 27:20]
  reg  vArrayWire_23_1; // @[Reg.scala 27:20]
  reg  vArrayWire_22_1; // @[Reg.scala 27:20]
  reg  vArrayWire_21_1; // @[Reg.scala 27:20]
  reg  vArrayWire_20_1; // @[Reg.scala 27:20]
  reg  vArrayWire_19_1; // @[Reg.scala 27:20]
  reg  vArrayWire_18_1; // @[Reg.scala 27:20]
  reg  vArrayWire_17_1; // @[Reg.scala 27:20]
  reg  vArrayWire_16_1; // @[Reg.scala 27:20]
  reg  vArrayWire_15_1; // @[Reg.scala 27:20]
  reg  vArrayWire_14_1; // @[Reg.scala 27:20]
  reg  vArrayWire_13_1; // @[Reg.scala 27:20]
  reg  vArrayWire_12_1; // @[Reg.scala 27:20]
  reg  vArrayWire_11_1; // @[Reg.scala 27:20]
  reg  vArrayWire_10_1; // @[Reg.scala 27:20]
  reg  vArrayWire_9_1; // @[Reg.scala 27:20]
  reg  vArrayWire_8_1; // @[Reg.scala 27:20]
  reg  vArrayWire_7_1; // @[Reg.scala 27:20]
  reg  vArrayWire_6_1; // @[Reg.scala 27:20]
  reg  vArrayWire_5_1; // @[Reg.scala 27:20]
  reg  vArrayWire_4_1; // @[Reg.scala 27:20]
  reg  vArrayWire_3_1; // @[Reg.scala 27:20]
  reg  vArrayWire_2_1; // @[Reg.scala 27:20]
  reg  vArrayWire_1_1; // @[Reg.scala 27:20]
  reg  vArrayWire_0_1; // @[Reg.scala 27:20]
  wire  _T_130_1 = _T_129 ? vArrayWire_1_1 : vArrayWire_0_1; // @[Mux.scala 80:57]
  wire  _T_132_1 = _T_131 ? vArrayWire_2_1 : _T_130_1; // @[Mux.scala 80:57]
  wire  _T_134_1 = _T_133 ? vArrayWire_3_1 : _T_132_1; // @[Mux.scala 80:57]
  wire  _T_136_1 = _T_135 ? vArrayWire_4_1 : _T_134_1; // @[Mux.scala 80:57]
  wire  _T_138_1 = _T_137 ? vArrayWire_5_1 : _T_136_1; // @[Mux.scala 80:57]
  wire  _T_140_1 = _T_139 ? vArrayWire_6_1 : _T_138_1; // @[Mux.scala 80:57]
  wire  _T_142_1 = _T_141 ? vArrayWire_7_1 : _T_140_1; // @[Mux.scala 80:57]
  wire  _T_144_1 = _T_143 ? vArrayWire_8_1 : _T_142_1; // @[Mux.scala 80:57]
  wire  _T_146_1 = _T_145 ? vArrayWire_9_1 : _T_144_1; // @[Mux.scala 80:57]
  wire  _T_148_1 = _T_147 ? vArrayWire_10_1 : _T_146_1; // @[Mux.scala 80:57]
  wire  _T_150_1 = _T_149 ? vArrayWire_11_1 : _T_148_1; // @[Mux.scala 80:57]
  wire  _T_152_1 = _T_151 ? vArrayWire_12_1 : _T_150_1; // @[Mux.scala 80:57]
  wire  _T_154_1 = _T_153 ? vArrayWire_13_1 : _T_152_1; // @[Mux.scala 80:57]
  wire  _T_156_1 = _T_155 ? vArrayWire_14_1 : _T_154_1; // @[Mux.scala 80:57]
  wire  _T_158_1 = _T_157 ? vArrayWire_15_1 : _T_156_1; // @[Mux.scala 80:57]
  wire  _T_160_1 = _T_159 ? vArrayWire_16_1 : _T_158_1; // @[Mux.scala 80:57]
  wire  _T_162_1 = _T_161 ? vArrayWire_17_1 : _T_160_1; // @[Mux.scala 80:57]
  wire  _T_164_1 = _T_163 ? vArrayWire_18_1 : _T_162_1; // @[Mux.scala 80:57]
  wire  _T_166_1 = _T_165 ? vArrayWire_19_1 : _T_164_1; // @[Mux.scala 80:57]
  wire  _T_168_1 = _T_167 ? vArrayWire_20_1 : _T_166_1; // @[Mux.scala 80:57]
  wire  _T_170_1 = _T_169 ? vArrayWire_21_1 : _T_168_1; // @[Mux.scala 80:57]
  wire  _T_172_1 = _T_171 ? vArrayWire_22_1 : _T_170_1; // @[Mux.scala 80:57]
  wire  _T_174_1 = _T_173 ? vArrayWire_23_1 : _T_172_1; // @[Mux.scala 80:57]
  wire  _T_176_1 = _T_175 ? vArrayWire_24_1 : _T_174_1; // @[Mux.scala 80:57]
  wire  _T_178_1 = _T_177 ? vArrayWire_25_1 : _T_176_1; // @[Mux.scala 80:57]
  wire  _T_180_1 = _T_179 ? vArrayWire_26_1 : _T_178_1; // @[Mux.scala 80:57]
  wire  _T_182_1 = _T_181 ? vArrayWire_27_1 : _T_180_1; // @[Mux.scala 80:57]
  wire  _T_184_1 = _T_183 ? vArrayWire_28_1 : _T_182_1; // @[Mux.scala 80:57]
  wire  _T_186_1 = _T_185 ? vArrayWire_29_1 : _T_184_1; // @[Mux.scala 80:57]
  wire  _T_188_1 = _T_187 ? vArrayWire_30_1 : _T_186_1; // @[Mux.scala 80:57]
  wire  _T_190_1 = _T_189 ? vArrayWire_31_1 : _T_188_1; // @[Mux.scala 80:57]
  wire  _T_192_1 = _T_191 ? vArrayWire_32_1 : _T_190_1; // @[Mux.scala 80:57]
  wire  _T_194_1 = _T_193 ? vArrayWire_33_1 : _T_192_1; // @[Mux.scala 80:57]
  wire  _T_196_1 = _T_195 ? vArrayWire_34_1 : _T_194_1; // @[Mux.scala 80:57]
  wire  _T_198_1 = _T_197 ? vArrayWire_35_1 : _T_196_1; // @[Mux.scala 80:57]
  wire  _T_200_1 = _T_199 ? vArrayWire_36_1 : _T_198_1; // @[Mux.scala 80:57]
  wire  _T_202_1 = _T_201 ? vArrayWire_37_1 : _T_200_1; // @[Mux.scala 80:57]
  wire  _T_204_1 = _T_203 ? vArrayWire_38_1 : _T_202_1; // @[Mux.scala 80:57]
  wire  _T_206_1 = _T_205 ? vArrayWire_39_1 : _T_204_1; // @[Mux.scala 80:57]
  wire  _T_208_1 = _T_207 ? vArrayWire_40_1 : _T_206_1; // @[Mux.scala 80:57]
  wire  _T_210_1 = _T_209 ? vArrayWire_41_1 : _T_208_1; // @[Mux.scala 80:57]
  wire  _T_212_1 = _T_211 ? vArrayWire_42_1 : _T_210_1; // @[Mux.scala 80:57]
  wire  _T_214_1 = _T_213 ? vArrayWire_43_1 : _T_212_1; // @[Mux.scala 80:57]
  wire  _T_216_1 = _T_215 ? vArrayWire_44_1 : _T_214_1; // @[Mux.scala 80:57]
  wire  _T_218_1 = _T_217 ? vArrayWire_45_1 : _T_216_1; // @[Mux.scala 80:57]
  wire  _T_220_1 = _T_219 ? vArrayWire_46_1 : _T_218_1; // @[Mux.scala 80:57]
  wire  _T_222_1 = _T_221 ? vArrayWire_47_1 : _T_220_1; // @[Mux.scala 80:57]
  wire  _T_224_1 = _T_223 ? vArrayWire_48_1 : _T_222_1; // @[Mux.scala 80:57]
  wire  _T_226_1 = _T_225 ? vArrayWire_49_1 : _T_224_1; // @[Mux.scala 80:57]
  wire  _T_228_1 = _T_227 ? vArrayWire_50_1 : _T_226_1; // @[Mux.scala 80:57]
  wire  _T_230_1 = _T_229 ? vArrayWire_51_1 : _T_228_1; // @[Mux.scala 80:57]
  wire  _T_232_1 = _T_231 ? vArrayWire_52_1 : _T_230_1; // @[Mux.scala 80:57]
  wire  _T_234_1 = _T_233 ? vArrayWire_53_1 : _T_232_1; // @[Mux.scala 80:57]
  wire  _T_236_1 = _T_235 ? vArrayWire_54_1 : _T_234_1; // @[Mux.scala 80:57]
  wire  _T_238_1 = _T_237 ? vArrayWire_55_1 : _T_236_1; // @[Mux.scala 80:57]
  wire  _T_240_1 = _T_239 ? vArrayWire_56_1 : _T_238_1; // @[Mux.scala 80:57]
  wire  _T_242_1 = _T_241 ? vArrayWire_57_1 : _T_240_1; // @[Mux.scala 80:57]
  wire  _T_244_1 = _T_243 ? vArrayWire_58_1 : _T_242_1; // @[Mux.scala 80:57]
  wire  _T_246_1 = _T_245 ? vArrayWire_59_1 : _T_244_1; // @[Mux.scala 80:57]
  wire  _T_248_1 = _T_247 ? vArrayWire_60_1 : _T_246_1; // @[Mux.scala 80:57]
  wire  _T_250_1 = _T_249 ? vArrayWire_61_1 : _T_248_1; // @[Mux.scala 80:57]
  wire  _T_252_1 = _T_251 ? vArrayWire_62_1 : _T_250_1; // @[Mux.scala 80:57]
  wire  vMuxOut_1 = _T_253 ? vArrayWire_63_1 : _T_252_1; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_1; // @[Reg.scala 27:20]
  wire [21:0] _T_5_1 = _T_129 ? tagArrayWire_1_1 : tagArrayWire_0_1; // @[Mux.scala 80:57]
  wire [21:0] _T_7_1 = _T_131 ? tagArrayWire_2_1 : _T_5_1; // @[Mux.scala 80:57]
  wire [21:0] _T_9_1 = _T_133 ? tagArrayWire_3_1 : _T_7_1; // @[Mux.scala 80:57]
  wire [21:0] _T_11_1 = _T_135 ? tagArrayWire_4_1 : _T_9_1; // @[Mux.scala 80:57]
  wire [21:0] _T_13_1 = _T_137 ? tagArrayWire_5_1 : _T_11_1; // @[Mux.scala 80:57]
  wire [21:0] _T_15_1 = _T_139 ? tagArrayWire_6_1 : _T_13_1; // @[Mux.scala 80:57]
  wire [21:0] _T_17_1 = _T_141 ? tagArrayWire_7_1 : _T_15_1; // @[Mux.scala 80:57]
  wire [21:0] _T_19_1 = _T_143 ? tagArrayWire_8_1 : _T_17_1; // @[Mux.scala 80:57]
  wire [21:0] _T_21_1 = _T_145 ? tagArrayWire_9_1 : _T_19_1; // @[Mux.scala 80:57]
  wire [21:0] _T_23_1 = _T_147 ? tagArrayWire_10_1 : _T_21_1; // @[Mux.scala 80:57]
  wire [21:0] _T_25_1 = _T_149 ? tagArrayWire_11_1 : _T_23_1; // @[Mux.scala 80:57]
  wire [21:0] _T_27_1 = _T_151 ? tagArrayWire_12_1 : _T_25_1; // @[Mux.scala 80:57]
  wire [21:0] _T_29_1 = _T_153 ? tagArrayWire_13_1 : _T_27_1; // @[Mux.scala 80:57]
  wire [21:0] _T_31_1 = _T_155 ? tagArrayWire_14_1 : _T_29_1; // @[Mux.scala 80:57]
  wire [21:0] _T_33_1 = _T_157 ? tagArrayWire_15_1 : _T_31_1; // @[Mux.scala 80:57]
  wire [21:0] _T_35_1 = _T_159 ? tagArrayWire_16_1 : _T_33_1; // @[Mux.scala 80:57]
  wire [21:0] _T_37_1 = _T_161 ? tagArrayWire_17_1 : _T_35_1; // @[Mux.scala 80:57]
  wire [21:0] _T_39_1 = _T_163 ? tagArrayWire_18_1 : _T_37_1; // @[Mux.scala 80:57]
  wire [21:0] _T_41_1 = _T_165 ? tagArrayWire_19_1 : _T_39_1; // @[Mux.scala 80:57]
  wire [21:0] _T_43_1 = _T_167 ? tagArrayWire_20_1 : _T_41_1; // @[Mux.scala 80:57]
  wire [21:0] _T_45_1 = _T_169 ? tagArrayWire_21_1 : _T_43_1; // @[Mux.scala 80:57]
  wire [21:0] _T_47_1 = _T_171 ? tagArrayWire_22_1 : _T_45_1; // @[Mux.scala 80:57]
  wire [21:0] _T_49_1 = _T_173 ? tagArrayWire_23_1 : _T_47_1; // @[Mux.scala 80:57]
  wire [21:0] _T_51_1 = _T_175 ? tagArrayWire_24_1 : _T_49_1; // @[Mux.scala 80:57]
  wire [21:0] _T_53_1 = _T_177 ? tagArrayWire_25_1 : _T_51_1; // @[Mux.scala 80:57]
  wire [21:0] _T_55_1 = _T_179 ? tagArrayWire_26_1 : _T_53_1; // @[Mux.scala 80:57]
  wire [21:0] _T_57_1 = _T_181 ? tagArrayWire_27_1 : _T_55_1; // @[Mux.scala 80:57]
  wire [21:0] _T_59_1 = _T_183 ? tagArrayWire_28_1 : _T_57_1; // @[Mux.scala 80:57]
  wire [21:0] _T_61_1 = _T_185 ? tagArrayWire_29_1 : _T_59_1; // @[Mux.scala 80:57]
  wire [21:0] _T_63_1 = _T_187 ? tagArrayWire_30_1 : _T_61_1; // @[Mux.scala 80:57]
  wire [21:0] _T_65_1 = _T_189 ? tagArrayWire_31_1 : _T_63_1; // @[Mux.scala 80:57]
  wire [21:0] _T_67_1 = _T_191 ? tagArrayWire_32_1 : _T_65_1; // @[Mux.scala 80:57]
  wire [21:0] _T_69_1 = _T_193 ? tagArrayWire_33_1 : _T_67_1; // @[Mux.scala 80:57]
  wire [21:0] _T_71_1 = _T_195 ? tagArrayWire_34_1 : _T_69_1; // @[Mux.scala 80:57]
  wire [21:0] _T_73_1 = _T_197 ? tagArrayWire_35_1 : _T_71_1; // @[Mux.scala 80:57]
  wire [21:0] _T_75_1 = _T_199 ? tagArrayWire_36_1 : _T_73_1; // @[Mux.scala 80:57]
  wire [21:0] _T_77_1 = _T_201 ? tagArrayWire_37_1 : _T_75_1; // @[Mux.scala 80:57]
  wire [21:0] _T_79_1 = _T_203 ? tagArrayWire_38_1 : _T_77_1; // @[Mux.scala 80:57]
  wire [21:0] _T_81_1 = _T_205 ? tagArrayWire_39_1 : _T_79_1; // @[Mux.scala 80:57]
  wire [21:0] _T_83_1 = _T_207 ? tagArrayWire_40_1 : _T_81_1; // @[Mux.scala 80:57]
  wire [21:0] _T_85_1 = _T_209 ? tagArrayWire_41_1 : _T_83_1; // @[Mux.scala 80:57]
  wire [21:0] _T_87_1 = _T_211 ? tagArrayWire_42_1 : _T_85_1; // @[Mux.scala 80:57]
  wire [21:0] _T_89_1 = _T_213 ? tagArrayWire_43_1 : _T_87_1; // @[Mux.scala 80:57]
  wire [21:0] _T_91_1 = _T_215 ? tagArrayWire_44_1 : _T_89_1; // @[Mux.scala 80:57]
  wire [21:0] _T_93_1 = _T_217 ? tagArrayWire_45_1 : _T_91_1; // @[Mux.scala 80:57]
  wire [21:0] _T_95_1 = _T_219 ? tagArrayWire_46_1 : _T_93_1; // @[Mux.scala 80:57]
  wire [21:0] _T_97_1 = _T_221 ? tagArrayWire_47_1 : _T_95_1; // @[Mux.scala 80:57]
  wire [21:0] _T_99_1 = _T_223 ? tagArrayWire_48_1 : _T_97_1; // @[Mux.scala 80:57]
  wire [21:0] _T_101_1 = _T_225 ? tagArrayWire_49_1 : _T_99_1; // @[Mux.scala 80:57]
  wire [21:0] _T_103_1 = _T_227 ? tagArrayWire_50_1 : _T_101_1; // @[Mux.scala 80:57]
  wire [21:0] _T_105_1 = _T_229 ? tagArrayWire_51_1 : _T_103_1; // @[Mux.scala 80:57]
  wire [21:0] _T_107_1 = _T_231 ? tagArrayWire_52_1 : _T_105_1; // @[Mux.scala 80:57]
  wire [21:0] _T_109_1 = _T_233 ? tagArrayWire_53_1 : _T_107_1; // @[Mux.scala 80:57]
  wire [21:0] _T_111_1 = _T_235 ? tagArrayWire_54_1 : _T_109_1; // @[Mux.scala 80:57]
  wire [21:0] _T_113_1 = _T_237 ? tagArrayWire_55_1 : _T_111_1; // @[Mux.scala 80:57]
  wire [21:0] _T_115_1 = _T_239 ? tagArrayWire_56_1 : _T_113_1; // @[Mux.scala 80:57]
  wire [21:0] _T_117_1 = _T_241 ? tagArrayWire_57_1 : _T_115_1; // @[Mux.scala 80:57]
  wire [21:0] _T_119_1 = _T_243 ? tagArrayWire_58_1 : _T_117_1; // @[Mux.scala 80:57]
  wire [21:0] _T_121_1 = _T_245 ? tagArrayWire_59_1 : _T_119_1; // @[Mux.scala 80:57]
  wire [21:0] _T_123_1 = _T_247 ? tagArrayWire_60_1 : _T_121_1; // @[Mux.scala 80:57]
  wire [21:0] _T_125_1 = _T_249 ? tagArrayWire_61_1 : _T_123_1; // @[Mux.scala 80:57]
  wire [21:0] _T_127_1 = _T_251 ? tagArrayWire_62_1 : _T_125_1; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_1 = _T_253 ? tagArrayWire_63_1 : _T_127_1; // @[Mux.scala 80:57]
  wire  _T_255 = tagMuxOut_1 == tag; // @[Cache.scala 72:76]
  wire  hitArray_1 = vMuxOut_1 & _T_255; // @[Cache.scala 72:60]
  wire  _T_259 = hitArray_0 | hitArray_1; // @[Cache.scala 73:49]
  reg  vArrayWire_63_2; // @[Reg.scala 27:20]
  reg  vArrayWire_62_2; // @[Reg.scala 27:20]
  reg  vArrayWire_61_2; // @[Reg.scala 27:20]
  reg  vArrayWire_60_2; // @[Reg.scala 27:20]
  reg  vArrayWire_59_2; // @[Reg.scala 27:20]
  reg  vArrayWire_58_2; // @[Reg.scala 27:20]
  reg  vArrayWire_57_2; // @[Reg.scala 27:20]
  reg  vArrayWire_56_2; // @[Reg.scala 27:20]
  reg  vArrayWire_55_2; // @[Reg.scala 27:20]
  reg  vArrayWire_54_2; // @[Reg.scala 27:20]
  reg  vArrayWire_53_2; // @[Reg.scala 27:20]
  reg  vArrayWire_52_2; // @[Reg.scala 27:20]
  reg  vArrayWire_51_2; // @[Reg.scala 27:20]
  reg  vArrayWire_50_2; // @[Reg.scala 27:20]
  reg  vArrayWire_49_2; // @[Reg.scala 27:20]
  reg  vArrayWire_48_2; // @[Reg.scala 27:20]
  reg  vArrayWire_47_2; // @[Reg.scala 27:20]
  reg  vArrayWire_46_2; // @[Reg.scala 27:20]
  reg  vArrayWire_45_2; // @[Reg.scala 27:20]
  reg  vArrayWire_44_2; // @[Reg.scala 27:20]
  reg  vArrayWire_43_2; // @[Reg.scala 27:20]
  reg  vArrayWire_42_2; // @[Reg.scala 27:20]
  reg  vArrayWire_41_2; // @[Reg.scala 27:20]
  reg  vArrayWire_40_2; // @[Reg.scala 27:20]
  reg  vArrayWire_39_2; // @[Reg.scala 27:20]
  reg  vArrayWire_38_2; // @[Reg.scala 27:20]
  reg  vArrayWire_37_2; // @[Reg.scala 27:20]
  reg  vArrayWire_36_2; // @[Reg.scala 27:20]
  reg  vArrayWire_35_2; // @[Reg.scala 27:20]
  reg  vArrayWire_34_2; // @[Reg.scala 27:20]
  reg  vArrayWire_33_2; // @[Reg.scala 27:20]
  reg  vArrayWire_32_2; // @[Reg.scala 27:20]
  reg  vArrayWire_31_2; // @[Reg.scala 27:20]
  reg  vArrayWire_30_2; // @[Reg.scala 27:20]
  reg  vArrayWire_29_2; // @[Reg.scala 27:20]
  reg  vArrayWire_28_2; // @[Reg.scala 27:20]
  reg  vArrayWire_27_2; // @[Reg.scala 27:20]
  reg  vArrayWire_26_2; // @[Reg.scala 27:20]
  reg  vArrayWire_25_2; // @[Reg.scala 27:20]
  reg  vArrayWire_24_2; // @[Reg.scala 27:20]
  reg  vArrayWire_23_2; // @[Reg.scala 27:20]
  reg  vArrayWire_22_2; // @[Reg.scala 27:20]
  reg  vArrayWire_21_2; // @[Reg.scala 27:20]
  reg  vArrayWire_20_2; // @[Reg.scala 27:20]
  reg  vArrayWire_19_2; // @[Reg.scala 27:20]
  reg  vArrayWire_18_2; // @[Reg.scala 27:20]
  reg  vArrayWire_17_2; // @[Reg.scala 27:20]
  reg  vArrayWire_16_2; // @[Reg.scala 27:20]
  reg  vArrayWire_15_2; // @[Reg.scala 27:20]
  reg  vArrayWire_14_2; // @[Reg.scala 27:20]
  reg  vArrayWire_13_2; // @[Reg.scala 27:20]
  reg  vArrayWire_12_2; // @[Reg.scala 27:20]
  reg  vArrayWire_11_2; // @[Reg.scala 27:20]
  reg  vArrayWire_10_2; // @[Reg.scala 27:20]
  reg  vArrayWire_9_2; // @[Reg.scala 27:20]
  reg  vArrayWire_8_2; // @[Reg.scala 27:20]
  reg  vArrayWire_7_2; // @[Reg.scala 27:20]
  reg  vArrayWire_6_2; // @[Reg.scala 27:20]
  reg  vArrayWire_5_2; // @[Reg.scala 27:20]
  reg  vArrayWire_4_2; // @[Reg.scala 27:20]
  reg  vArrayWire_3_2; // @[Reg.scala 27:20]
  reg  vArrayWire_2_2; // @[Reg.scala 27:20]
  reg  vArrayWire_1_2; // @[Reg.scala 27:20]
  reg  vArrayWire_0_2; // @[Reg.scala 27:20]
  wire  _T_130_2 = _T_129 ? vArrayWire_1_2 : vArrayWire_0_2; // @[Mux.scala 80:57]
  wire  _T_132_2 = _T_131 ? vArrayWire_2_2 : _T_130_2; // @[Mux.scala 80:57]
  wire  _T_134_2 = _T_133 ? vArrayWire_3_2 : _T_132_2; // @[Mux.scala 80:57]
  wire  _T_136_2 = _T_135 ? vArrayWire_4_2 : _T_134_2; // @[Mux.scala 80:57]
  wire  _T_138_2 = _T_137 ? vArrayWire_5_2 : _T_136_2; // @[Mux.scala 80:57]
  wire  _T_140_2 = _T_139 ? vArrayWire_6_2 : _T_138_2; // @[Mux.scala 80:57]
  wire  _T_142_2 = _T_141 ? vArrayWire_7_2 : _T_140_2; // @[Mux.scala 80:57]
  wire  _T_144_2 = _T_143 ? vArrayWire_8_2 : _T_142_2; // @[Mux.scala 80:57]
  wire  _T_146_2 = _T_145 ? vArrayWire_9_2 : _T_144_2; // @[Mux.scala 80:57]
  wire  _T_148_2 = _T_147 ? vArrayWire_10_2 : _T_146_2; // @[Mux.scala 80:57]
  wire  _T_150_2 = _T_149 ? vArrayWire_11_2 : _T_148_2; // @[Mux.scala 80:57]
  wire  _T_152_2 = _T_151 ? vArrayWire_12_2 : _T_150_2; // @[Mux.scala 80:57]
  wire  _T_154_2 = _T_153 ? vArrayWire_13_2 : _T_152_2; // @[Mux.scala 80:57]
  wire  _T_156_2 = _T_155 ? vArrayWire_14_2 : _T_154_2; // @[Mux.scala 80:57]
  wire  _T_158_2 = _T_157 ? vArrayWire_15_2 : _T_156_2; // @[Mux.scala 80:57]
  wire  _T_160_2 = _T_159 ? vArrayWire_16_2 : _T_158_2; // @[Mux.scala 80:57]
  wire  _T_162_2 = _T_161 ? vArrayWire_17_2 : _T_160_2; // @[Mux.scala 80:57]
  wire  _T_164_2 = _T_163 ? vArrayWire_18_2 : _T_162_2; // @[Mux.scala 80:57]
  wire  _T_166_2 = _T_165 ? vArrayWire_19_2 : _T_164_2; // @[Mux.scala 80:57]
  wire  _T_168_2 = _T_167 ? vArrayWire_20_2 : _T_166_2; // @[Mux.scala 80:57]
  wire  _T_170_2 = _T_169 ? vArrayWire_21_2 : _T_168_2; // @[Mux.scala 80:57]
  wire  _T_172_2 = _T_171 ? vArrayWire_22_2 : _T_170_2; // @[Mux.scala 80:57]
  wire  _T_174_2 = _T_173 ? vArrayWire_23_2 : _T_172_2; // @[Mux.scala 80:57]
  wire  _T_176_2 = _T_175 ? vArrayWire_24_2 : _T_174_2; // @[Mux.scala 80:57]
  wire  _T_178_2 = _T_177 ? vArrayWire_25_2 : _T_176_2; // @[Mux.scala 80:57]
  wire  _T_180_2 = _T_179 ? vArrayWire_26_2 : _T_178_2; // @[Mux.scala 80:57]
  wire  _T_182_2 = _T_181 ? vArrayWire_27_2 : _T_180_2; // @[Mux.scala 80:57]
  wire  _T_184_2 = _T_183 ? vArrayWire_28_2 : _T_182_2; // @[Mux.scala 80:57]
  wire  _T_186_2 = _T_185 ? vArrayWire_29_2 : _T_184_2; // @[Mux.scala 80:57]
  wire  _T_188_2 = _T_187 ? vArrayWire_30_2 : _T_186_2; // @[Mux.scala 80:57]
  wire  _T_190_2 = _T_189 ? vArrayWire_31_2 : _T_188_2; // @[Mux.scala 80:57]
  wire  _T_192_2 = _T_191 ? vArrayWire_32_2 : _T_190_2; // @[Mux.scala 80:57]
  wire  _T_194_2 = _T_193 ? vArrayWire_33_2 : _T_192_2; // @[Mux.scala 80:57]
  wire  _T_196_2 = _T_195 ? vArrayWire_34_2 : _T_194_2; // @[Mux.scala 80:57]
  wire  _T_198_2 = _T_197 ? vArrayWire_35_2 : _T_196_2; // @[Mux.scala 80:57]
  wire  _T_200_2 = _T_199 ? vArrayWire_36_2 : _T_198_2; // @[Mux.scala 80:57]
  wire  _T_202_2 = _T_201 ? vArrayWire_37_2 : _T_200_2; // @[Mux.scala 80:57]
  wire  _T_204_2 = _T_203 ? vArrayWire_38_2 : _T_202_2; // @[Mux.scala 80:57]
  wire  _T_206_2 = _T_205 ? vArrayWire_39_2 : _T_204_2; // @[Mux.scala 80:57]
  wire  _T_208_2 = _T_207 ? vArrayWire_40_2 : _T_206_2; // @[Mux.scala 80:57]
  wire  _T_210_2 = _T_209 ? vArrayWire_41_2 : _T_208_2; // @[Mux.scala 80:57]
  wire  _T_212_2 = _T_211 ? vArrayWire_42_2 : _T_210_2; // @[Mux.scala 80:57]
  wire  _T_214_2 = _T_213 ? vArrayWire_43_2 : _T_212_2; // @[Mux.scala 80:57]
  wire  _T_216_2 = _T_215 ? vArrayWire_44_2 : _T_214_2; // @[Mux.scala 80:57]
  wire  _T_218_2 = _T_217 ? vArrayWire_45_2 : _T_216_2; // @[Mux.scala 80:57]
  wire  _T_220_2 = _T_219 ? vArrayWire_46_2 : _T_218_2; // @[Mux.scala 80:57]
  wire  _T_222_2 = _T_221 ? vArrayWire_47_2 : _T_220_2; // @[Mux.scala 80:57]
  wire  _T_224_2 = _T_223 ? vArrayWire_48_2 : _T_222_2; // @[Mux.scala 80:57]
  wire  _T_226_2 = _T_225 ? vArrayWire_49_2 : _T_224_2; // @[Mux.scala 80:57]
  wire  _T_228_2 = _T_227 ? vArrayWire_50_2 : _T_226_2; // @[Mux.scala 80:57]
  wire  _T_230_2 = _T_229 ? vArrayWire_51_2 : _T_228_2; // @[Mux.scala 80:57]
  wire  _T_232_2 = _T_231 ? vArrayWire_52_2 : _T_230_2; // @[Mux.scala 80:57]
  wire  _T_234_2 = _T_233 ? vArrayWire_53_2 : _T_232_2; // @[Mux.scala 80:57]
  wire  _T_236_2 = _T_235 ? vArrayWire_54_2 : _T_234_2; // @[Mux.scala 80:57]
  wire  _T_238_2 = _T_237 ? vArrayWire_55_2 : _T_236_2; // @[Mux.scala 80:57]
  wire  _T_240_2 = _T_239 ? vArrayWire_56_2 : _T_238_2; // @[Mux.scala 80:57]
  wire  _T_242_2 = _T_241 ? vArrayWire_57_2 : _T_240_2; // @[Mux.scala 80:57]
  wire  _T_244_2 = _T_243 ? vArrayWire_58_2 : _T_242_2; // @[Mux.scala 80:57]
  wire  _T_246_2 = _T_245 ? vArrayWire_59_2 : _T_244_2; // @[Mux.scala 80:57]
  wire  _T_248_2 = _T_247 ? vArrayWire_60_2 : _T_246_2; // @[Mux.scala 80:57]
  wire  _T_250_2 = _T_249 ? vArrayWire_61_2 : _T_248_2; // @[Mux.scala 80:57]
  wire  _T_252_2 = _T_251 ? vArrayWire_62_2 : _T_250_2; // @[Mux.scala 80:57]
  wire  vMuxOut_2 = _T_253 ? vArrayWire_63_2 : _T_252_2; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_2; // @[Reg.scala 27:20]
  wire [21:0] _T_5_2 = _T_129 ? tagArrayWire_1_2 : tagArrayWire_0_2; // @[Mux.scala 80:57]
  wire [21:0] _T_7_2 = _T_131 ? tagArrayWire_2_2 : _T_5_2; // @[Mux.scala 80:57]
  wire [21:0] _T_9_2 = _T_133 ? tagArrayWire_3_2 : _T_7_2; // @[Mux.scala 80:57]
  wire [21:0] _T_11_2 = _T_135 ? tagArrayWire_4_2 : _T_9_2; // @[Mux.scala 80:57]
  wire [21:0] _T_13_2 = _T_137 ? tagArrayWire_5_2 : _T_11_2; // @[Mux.scala 80:57]
  wire [21:0] _T_15_2 = _T_139 ? tagArrayWire_6_2 : _T_13_2; // @[Mux.scala 80:57]
  wire [21:0] _T_17_2 = _T_141 ? tagArrayWire_7_2 : _T_15_2; // @[Mux.scala 80:57]
  wire [21:0] _T_19_2 = _T_143 ? tagArrayWire_8_2 : _T_17_2; // @[Mux.scala 80:57]
  wire [21:0] _T_21_2 = _T_145 ? tagArrayWire_9_2 : _T_19_2; // @[Mux.scala 80:57]
  wire [21:0] _T_23_2 = _T_147 ? tagArrayWire_10_2 : _T_21_2; // @[Mux.scala 80:57]
  wire [21:0] _T_25_2 = _T_149 ? tagArrayWire_11_2 : _T_23_2; // @[Mux.scala 80:57]
  wire [21:0] _T_27_2 = _T_151 ? tagArrayWire_12_2 : _T_25_2; // @[Mux.scala 80:57]
  wire [21:0] _T_29_2 = _T_153 ? tagArrayWire_13_2 : _T_27_2; // @[Mux.scala 80:57]
  wire [21:0] _T_31_2 = _T_155 ? tagArrayWire_14_2 : _T_29_2; // @[Mux.scala 80:57]
  wire [21:0] _T_33_2 = _T_157 ? tagArrayWire_15_2 : _T_31_2; // @[Mux.scala 80:57]
  wire [21:0] _T_35_2 = _T_159 ? tagArrayWire_16_2 : _T_33_2; // @[Mux.scala 80:57]
  wire [21:0] _T_37_2 = _T_161 ? tagArrayWire_17_2 : _T_35_2; // @[Mux.scala 80:57]
  wire [21:0] _T_39_2 = _T_163 ? tagArrayWire_18_2 : _T_37_2; // @[Mux.scala 80:57]
  wire [21:0] _T_41_2 = _T_165 ? tagArrayWire_19_2 : _T_39_2; // @[Mux.scala 80:57]
  wire [21:0] _T_43_2 = _T_167 ? tagArrayWire_20_2 : _T_41_2; // @[Mux.scala 80:57]
  wire [21:0] _T_45_2 = _T_169 ? tagArrayWire_21_2 : _T_43_2; // @[Mux.scala 80:57]
  wire [21:0] _T_47_2 = _T_171 ? tagArrayWire_22_2 : _T_45_2; // @[Mux.scala 80:57]
  wire [21:0] _T_49_2 = _T_173 ? tagArrayWire_23_2 : _T_47_2; // @[Mux.scala 80:57]
  wire [21:0] _T_51_2 = _T_175 ? tagArrayWire_24_2 : _T_49_2; // @[Mux.scala 80:57]
  wire [21:0] _T_53_2 = _T_177 ? tagArrayWire_25_2 : _T_51_2; // @[Mux.scala 80:57]
  wire [21:0] _T_55_2 = _T_179 ? tagArrayWire_26_2 : _T_53_2; // @[Mux.scala 80:57]
  wire [21:0] _T_57_2 = _T_181 ? tagArrayWire_27_2 : _T_55_2; // @[Mux.scala 80:57]
  wire [21:0] _T_59_2 = _T_183 ? tagArrayWire_28_2 : _T_57_2; // @[Mux.scala 80:57]
  wire [21:0] _T_61_2 = _T_185 ? tagArrayWire_29_2 : _T_59_2; // @[Mux.scala 80:57]
  wire [21:0] _T_63_2 = _T_187 ? tagArrayWire_30_2 : _T_61_2; // @[Mux.scala 80:57]
  wire [21:0] _T_65_2 = _T_189 ? tagArrayWire_31_2 : _T_63_2; // @[Mux.scala 80:57]
  wire [21:0] _T_67_2 = _T_191 ? tagArrayWire_32_2 : _T_65_2; // @[Mux.scala 80:57]
  wire [21:0] _T_69_2 = _T_193 ? tagArrayWire_33_2 : _T_67_2; // @[Mux.scala 80:57]
  wire [21:0] _T_71_2 = _T_195 ? tagArrayWire_34_2 : _T_69_2; // @[Mux.scala 80:57]
  wire [21:0] _T_73_2 = _T_197 ? tagArrayWire_35_2 : _T_71_2; // @[Mux.scala 80:57]
  wire [21:0] _T_75_2 = _T_199 ? tagArrayWire_36_2 : _T_73_2; // @[Mux.scala 80:57]
  wire [21:0] _T_77_2 = _T_201 ? tagArrayWire_37_2 : _T_75_2; // @[Mux.scala 80:57]
  wire [21:0] _T_79_2 = _T_203 ? tagArrayWire_38_2 : _T_77_2; // @[Mux.scala 80:57]
  wire [21:0] _T_81_2 = _T_205 ? tagArrayWire_39_2 : _T_79_2; // @[Mux.scala 80:57]
  wire [21:0] _T_83_2 = _T_207 ? tagArrayWire_40_2 : _T_81_2; // @[Mux.scala 80:57]
  wire [21:0] _T_85_2 = _T_209 ? tagArrayWire_41_2 : _T_83_2; // @[Mux.scala 80:57]
  wire [21:0] _T_87_2 = _T_211 ? tagArrayWire_42_2 : _T_85_2; // @[Mux.scala 80:57]
  wire [21:0] _T_89_2 = _T_213 ? tagArrayWire_43_2 : _T_87_2; // @[Mux.scala 80:57]
  wire [21:0] _T_91_2 = _T_215 ? tagArrayWire_44_2 : _T_89_2; // @[Mux.scala 80:57]
  wire [21:0] _T_93_2 = _T_217 ? tagArrayWire_45_2 : _T_91_2; // @[Mux.scala 80:57]
  wire [21:0] _T_95_2 = _T_219 ? tagArrayWire_46_2 : _T_93_2; // @[Mux.scala 80:57]
  wire [21:0] _T_97_2 = _T_221 ? tagArrayWire_47_2 : _T_95_2; // @[Mux.scala 80:57]
  wire [21:0] _T_99_2 = _T_223 ? tagArrayWire_48_2 : _T_97_2; // @[Mux.scala 80:57]
  wire [21:0] _T_101_2 = _T_225 ? tagArrayWire_49_2 : _T_99_2; // @[Mux.scala 80:57]
  wire [21:0] _T_103_2 = _T_227 ? tagArrayWire_50_2 : _T_101_2; // @[Mux.scala 80:57]
  wire [21:0] _T_105_2 = _T_229 ? tagArrayWire_51_2 : _T_103_2; // @[Mux.scala 80:57]
  wire [21:0] _T_107_2 = _T_231 ? tagArrayWire_52_2 : _T_105_2; // @[Mux.scala 80:57]
  wire [21:0] _T_109_2 = _T_233 ? tagArrayWire_53_2 : _T_107_2; // @[Mux.scala 80:57]
  wire [21:0] _T_111_2 = _T_235 ? tagArrayWire_54_2 : _T_109_2; // @[Mux.scala 80:57]
  wire [21:0] _T_113_2 = _T_237 ? tagArrayWire_55_2 : _T_111_2; // @[Mux.scala 80:57]
  wire [21:0] _T_115_2 = _T_239 ? tagArrayWire_56_2 : _T_113_2; // @[Mux.scala 80:57]
  wire [21:0] _T_117_2 = _T_241 ? tagArrayWire_57_2 : _T_115_2; // @[Mux.scala 80:57]
  wire [21:0] _T_119_2 = _T_243 ? tagArrayWire_58_2 : _T_117_2; // @[Mux.scala 80:57]
  wire [21:0] _T_121_2 = _T_245 ? tagArrayWire_59_2 : _T_119_2; // @[Mux.scala 80:57]
  wire [21:0] _T_123_2 = _T_247 ? tagArrayWire_60_2 : _T_121_2; // @[Mux.scala 80:57]
  wire [21:0] _T_125_2 = _T_249 ? tagArrayWire_61_2 : _T_123_2; // @[Mux.scala 80:57]
  wire [21:0] _T_127_2 = _T_251 ? tagArrayWire_62_2 : _T_125_2; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_2 = _T_253 ? tagArrayWire_63_2 : _T_127_2; // @[Mux.scala 80:57]
  wire  _T_256 = tagMuxOut_2 == tag; // @[Cache.scala 72:76]
  wire  hitArray_2 = vMuxOut_2 & _T_256; // @[Cache.scala 72:60]
  wire  _T_260 = _T_259 | hitArray_2; // @[Cache.scala 73:49]
  reg  vArrayWire_63_3; // @[Reg.scala 27:20]
  reg  vArrayWire_62_3; // @[Reg.scala 27:20]
  reg  vArrayWire_61_3; // @[Reg.scala 27:20]
  reg  vArrayWire_60_3; // @[Reg.scala 27:20]
  reg  vArrayWire_59_3; // @[Reg.scala 27:20]
  reg  vArrayWire_58_3; // @[Reg.scala 27:20]
  reg  vArrayWire_57_3; // @[Reg.scala 27:20]
  reg  vArrayWire_56_3; // @[Reg.scala 27:20]
  reg  vArrayWire_55_3; // @[Reg.scala 27:20]
  reg  vArrayWire_54_3; // @[Reg.scala 27:20]
  reg  vArrayWire_53_3; // @[Reg.scala 27:20]
  reg  vArrayWire_52_3; // @[Reg.scala 27:20]
  reg  vArrayWire_51_3; // @[Reg.scala 27:20]
  reg  vArrayWire_50_3; // @[Reg.scala 27:20]
  reg  vArrayWire_49_3; // @[Reg.scala 27:20]
  reg  vArrayWire_48_3; // @[Reg.scala 27:20]
  reg  vArrayWire_47_3; // @[Reg.scala 27:20]
  reg  vArrayWire_46_3; // @[Reg.scala 27:20]
  reg  vArrayWire_45_3; // @[Reg.scala 27:20]
  reg  vArrayWire_44_3; // @[Reg.scala 27:20]
  reg  vArrayWire_43_3; // @[Reg.scala 27:20]
  reg  vArrayWire_42_3; // @[Reg.scala 27:20]
  reg  vArrayWire_41_3; // @[Reg.scala 27:20]
  reg  vArrayWire_40_3; // @[Reg.scala 27:20]
  reg  vArrayWire_39_3; // @[Reg.scala 27:20]
  reg  vArrayWire_38_3; // @[Reg.scala 27:20]
  reg  vArrayWire_37_3; // @[Reg.scala 27:20]
  reg  vArrayWire_36_3; // @[Reg.scala 27:20]
  reg  vArrayWire_35_3; // @[Reg.scala 27:20]
  reg  vArrayWire_34_3; // @[Reg.scala 27:20]
  reg  vArrayWire_33_3; // @[Reg.scala 27:20]
  reg  vArrayWire_32_3; // @[Reg.scala 27:20]
  reg  vArrayWire_31_3; // @[Reg.scala 27:20]
  reg  vArrayWire_30_3; // @[Reg.scala 27:20]
  reg  vArrayWire_29_3; // @[Reg.scala 27:20]
  reg  vArrayWire_28_3; // @[Reg.scala 27:20]
  reg  vArrayWire_27_3; // @[Reg.scala 27:20]
  reg  vArrayWire_26_3; // @[Reg.scala 27:20]
  reg  vArrayWire_25_3; // @[Reg.scala 27:20]
  reg  vArrayWire_24_3; // @[Reg.scala 27:20]
  reg  vArrayWire_23_3; // @[Reg.scala 27:20]
  reg  vArrayWire_22_3; // @[Reg.scala 27:20]
  reg  vArrayWire_21_3; // @[Reg.scala 27:20]
  reg  vArrayWire_20_3; // @[Reg.scala 27:20]
  reg  vArrayWire_19_3; // @[Reg.scala 27:20]
  reg  vArrayWire_18_3; // @[Reg.scala 27:20]
  reg  vArrayWire_17_3; // @[Reg.scala 27:20]
  reg  vArrayWire_16_3; // @[Reg.scala 27:20]
  reg  vArrayWire_15_3; // @[Reg.scala 27:20]
  reg  vArrayWire_14_3; // @[Reg.scala 27:20]
  reg  vArrayWire_13_3; // @[Reg.scala 27:20]
  reg  vArrayWire_12_3; // @[Reg.scala 27:20]
  reg  vArrayWire_11_3; // @[Reg.scala 27:20]
  reg  vArrayWire_10_3; // @[Reg.scala 27:20]
  reg  vArrayWire_9_3; // @[Reg.scala 27:20]
  reg  vArrayWire_8_3; // @[Reg.scala 27:20]
  reg  vArrayWire_7_3; // @[Reg.scala 27:20]
  reg  vArrayWire_6_3; // @[Reg.scala 27:20]
  reg  vArrayWire_5_3; // @[Reg.scala 27:20]
  reg  vArrayWire_4_3; // @[Reg.scala 27:20]
  reg  vArrayWire_3_3; // @[Reg.scala 27:20]
  reg  vArrayWire_2_3; // @[Reg.scala 27:20]
  reg  vArrayWire_1_3; // @[Reg.scala 27:20]
  reg  vArrayWire_0_3; // @[Reg.scala 27:20]
  wire  _T_130_3 = _T_129 ? vArrayWire_1_3 : vArrayWire_0_3; // @[Mux.scala 80:57]
  wire  _T_132_3 = _T_131 ? vArrayWire_2_3 : _T_130_3; // @[Mux.scala 80:57]
  wire  _T_134_3 = _T_133 ? vArrayWire_3_3 : _T_132_3; // @[Mux.scala 80:57]
  wire  _T_136_3 = _T_135 ? vArrayWire_4_3 : _T_134_3; // @[Mux.scala 80:57]
  wire  _T_138_3 = _T_137 ? vArrayWire_5_3 : _T_136_3; // @[Mux.scala 80:57]
  wire  _T_140_3 = _T_139 ? vArrayWire_6_3 : _T_138_3; // @[Mux.scala 80:57]
  wire  _T_142_3 = _T_141 ? vArrayWire_7_3 : _T_140_3; // @[Mux.scala 80:57]
  wire  _T_144_3 = _T_143 ? vArrayWire_8_3 : _T_142_3; // @[Mux.scala 80:57]
  wire  _T_146_3 = _T_145 ? vArrayWire_9_3 : _T_144_3; // @[Mux.scala 80:57]
  wire  _T_148_3 = _T_147 ? vArrayWire_10_3 : _T_146_3; // @[Mux.scala 80:57]
  wire  _T_150_3 = _T_149 ? vArrayWire_11_3 : _T_148_3; // @[Mux.scala 80:57]
  wire  _T_152_3 = _T_151 ? vArrayWire_12_3 : _T_150_3; // @[Mux.scala 80:57]
  wire  _T_154_3 = _T_153 ? vArrayWire_13_3 : _T_152_3; // @[Mux.scala 80:57]
  wire  _T_156_3 = _T_155 ? vArrayWire_14_3 : _T_154_3; // @[Mux.scala 80:57]
  wire  _T_158_3 = _T_157 ? vArrayWire_15_3 : _T_156_3; // @[Mux.scala 80:57]
  wire  _T_160_3 = _T_159 ? vArrayWire_16_3 : _T_158_3; // @[Mux.scala 80:57]
  wire  _T_162_3 = _T_161 ? vArrayWire_17_3 : _T_160_3; // @[Mux.scala 80:57]
  wire  _T_164_3 = _T_163 ? vArrayWire_18_3 : _T_162_3; // @[Mux.scala 80:57]
  wire  _T_166_3 = _T_165 ? vArrayWire_19_3 : _T_164_3; // @[Mux.scala 80:57]
  wire  _T_168_3 = _T_167 ? vArrayWire_20_3 : _T_166_3; // @[Mux.scala 80:57]
  wire  _T_170_3 = _T_169 ? vArrayWire_21_3 : _T_168_3; // @[Mux.scala 80:57]
  wire  _T_172_3 = _T_171 ? vArrayWire_22_3 : _T_170_3; // @[Mux.scala 80:57]
  wire  _T_174_3 = _T_173 ? vArrayWire_23_3 : _T_172_3; // @[Mux.scala 80:57]
  wire  _T_176_3 = _T_175 ? vArrayWire_24_3 : _T_174_3; // @[Mux.scala 80:57]
  wire  _T_178_3 = _T_177 ? vArrayWire_25_3 : _T_176_3; // @[Mux.scala 80:57]
  wire  _T_180_3 = _T_179 ? vArrayWire_26_3 : _T_178_3; // @[Mux.scala 80:57]
  wire  _T_182_3 = _T_181 ? vArrayWire_27_3 : _T_180_3; // @[Mux.scala 80:57]
  wire  _T_184_3 = _T_183 ? vArrayWire_28_3 : _T_182_3; // @[Mux.scala 80:57]
  wire  _T_186_3 = _T_185 ? vArrayWire_29_3 : _T_184_3; // @[Mux.scala 80:57]
  wire  _T_188_3 = _T_187 ? vArrayWire_30_3 : _T_186_3; // @[Mux.scala 80:57]
  wire  _T_190_3 = _T_189 ? vArrayWire_31_3 : _T_188_3; // @[Mux.scala 80:57]
  wire  _T_192_3 = _T_191 ? vArrayWire_32_3 : _T_190_3; // @[Mux.scala 80:57]
  wire  _T_194_3 = _T_193 ? vArrayWire_33_3 : _T_192_3; // @[Mux.scala 80:57]
  wire  _T_196_3 = _T_195 ? vArrayWire_34_3 : _T_194_3; // @[Mux.scala 80:57]
  wire  _T_198_3 = _T_197 ? vArrayWire_35_3 : _T_196_3; // @[Mux.scala 80:57]
  wire  _T_200_3 = _T_199 ? vArrayWire_36_3 : _T_198_3; // @[Mux.scala 80:57]
  wire  _T_202_3 = _T_201 ? vArrayWire_37_3 : _T_200_3; // @[Mux.scala 80:57]
  wire  _T_204_3 = _T_203 ? vArrayWire_38_3 : _T_202_3; // @[Mux.scala 80:57]
  wire  _T_206_3 = _T_205 ? vArrayWire_39_3 : _T_204_3; // @[Mux.scala 80:57]
  wire  _T_208_3 = _T_207 ? vArrayWire_40_3 : _T_206_3; // @[Mux.scala 80:57]
  wire  _T_210_3 = _T_209 ? vArrayWire_41_3 : _T_208_3; // @[Mux.scala 80:57]
  wire  _T_212_3 = _T_211 ? vArrayWire_42_3 : _T_210_3; // @[Mux.scala 80:57]
  wire  _T_214_3 = _T_213 ? vArrayWire_43_3 : _T_212_3; // @[Mux.scala 80:57]
  wire  _T_216_3 = _T_215 ? vArrayWire_44_3 : _T_214_3; // @[Mux.scala 80:57]
  wire  _T_218_3 = _T_217 ? vArrayWire_45_3 : _T_216_3; // @[Mux.scala 80:57]
  wire  _T_220_3 = _T_219 ? vArrayWire_46_3 : _T_218_3; // @[Mux.scala 80:57]
  wire  _T_222_3 = _T_221 ? vArrayWire_47_3 : _T_220_3; // @[Mux.scala 80:57]
  wire  _T_224_3 = _T_223 ? vArrayWire_48_3 : _T_222_3; // @[Mux.scala 80:57]
  wire  _T_226_3 = _T_225 ? vArrayWire_49_3 : _T_224_3; // @[Mux.scala 80:57]
  wire  _T_228_3 = _T_227 ? vArrayWire_50_3 : _T_226_3; // @[Mux.scala 80:57]
  wire  _T_230_3 = _T_229 ? vArrayWire_51_3 : _T_228_3; // @[Mux.scala 80:57]
  wire  _T_232_3 = _T_231 ? vArrayWire_52_3 : _T_230_3; // @[Mux.scala 80:57]
  wire  _T_234_3 = _T_233 ? vArrayWire_53_3 : _T_232_3; // @[Mux.scala 80:57]
  wire  _T_236_3 = _T_235 ? vArrayWire_54_3 : _T_234_3; // @[Mux.scala 80:57]
  wire  _T_238_3 = _T_237 ? vArrayWire_55_3 : _T_236_3; // @[Mux.scala 80:57]
  wire  _T_240_3 = _T_239 ? vArrayWire_56_3 : _T_238_3; // @[Mux.scala 80:57]
  wire  _T_242_3 = _T_241 ? vArrayWire_57_3 : _T_240_3; // @[Mux.scala 80:57]
  wire  _T_244_3 = _T_243 ? vArrayWire_58_3 : _T_242_3; // @[Mux.scala 80:57]
  wire  _T_246_3 = _T_245 ? vArrayWire_59_3 : _T_244_3; // @[Mux.scala 80:57]
  wire  _T_248_3 = _T_247 ? vArrayWire_60_3 : _T_246_3; // @[Mux.scala 80:57]
  wire  _T_250_3 = _T_249 ? vArrayWire_61_3 : _T_248_3; // @[Mux.scala 80:57]
  wire  _T_252_3 = _T_251 ? vArrayWire_62_3 : _T_250_3; // @[Mux.scala 80:57]
  wire  vMuxOut_3 = _T_253 ? vArrayWire_63_3 : _T_252_3; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_3; // @[Reg.scala 27:20]
  wire [21:0] _T_5_3 = _T_129 ? tagArrayWire_1_3 : tagArrayWire_0_3; // @[Mux.scala 80:57]
  wire [21:0] _T_7_3 = _T_131 ? tagArrayWire_2_3 : _T_5_3; // @[Mux.scala 80:57]
  wire [21:0] _T_9_3 = _T_133 ? tagArrayWire_3_3 : _T_7_3; // @[Mux.scala 80:57]
  wire [21:0] _T_11_3 = _T_135 ? tagArrayWire_4_3 : _T_9_3; // @[Mux.scala 80:57]
  wire [21:0] _T_13_3 = _T_137 ? tagArrayWire_5_3 : _T_11_3; // @[Mux.scala 80:57]
  wire [21:0] _T_15_3 = _T_139 ? tagArrayWire_6_3 : _T_13_3; // @[Mux.scala 80:57]
  wire [21:0] _T_17_3 = _T_141 ? tagArrayWire_7_3 : _T_15_3; // @[Mux.scala 80:57]
  wire [21:0] _T_19_3 = _T_143 ? tagArrayWire_8_3 : _T_17_3; // @[Mux.scala 80:57]
  wire [21:0] _T_21_3 = _T_145 ? tagArrayWire_9_3 : _T_19_3; // @[Mux.scala 80:57]
  wire [21:0] _T_23_3 = _T_147 ? tagArrayWire_10_3 : _T_21_3; // @[Mux.scala 80:57]
  wire [21:0] _T_25_3 = _T_149 ? tagArrayWire_11_3 : _T_23_3; // @[Mux.scala 80:57]
  wire [21:0] _T_27_3 = _T_151 ? tagArrayWire_12_3 : _T_25_3; // @[Mux.scala 80:57]
  wire [21:0] _T_29_3 = _T_153 ? tagArrayWire_13_3 : _T_27_3; // @[Mux.scala 80:57]
  wire [21:0] _T_31_3 = _T_155 ? tagArrayWire_14_3 : _T_29_3; // @[Mux.scala 80:57]
  wire [21:0] _T_33_3 = _T_157 ? tagArrayWire_15_3 : _T_31_3; // @[Mux.scala 80:57]
  wire [21:0] _T_35_3 = _T_159 ? tagArrayWire_16_3 : _T_33_3; // @[Mux.scala 80:57]
  wire [21:0] _T_37_3 = _T_161 ? tagArrayWire_17_3 : _T_35_3; // @[Mux.scala 80:57]
  wire [21:0] _T_39_3 = _T_163 ? tagArrayWire_18_3 : _T_37_3; // @[Mux.scala 80:57]
  wire [21:0] _T_41_3 = _T_165 ? tagArrayWire_19_3 : _T_39_3; // @[Mux.scala 80:57]
  wire [21:0] _T_43_3 = _T_167 ? tagArrayWire_20_3 : _T_41_3; // @[Mux.scala 80:57]
  wire [21:0] _T_45_3 = _T_169 ? tagArrayWire_21_3 : _T_43_3; // @[Mux.scala 80:57]
  wire [21:0] _T_47_3 = _T_171 ? tagArrayWire_22_3 : _T_45_3; // @[Mux.scala 80:57]
  wire [21:0] _T_49_3 = _T_173 ? tagArrayWire_23_3 : _T_47_3; // @[Mux.scala 80:57]
  wire [21:0] _T_51_3 = _T_175 ? tagArrayWire_24_3 : _T_49_3; // @[Mux.scala 80:57]
  wire [21:0] _T_53_3 = _T_177 ? tagArrayWire_25_3 : _T_51_3; // @[Mux.scala 80:57]
  wire [21:0] _T_55_3 = _T_179 ? tagArrayWire_26_3 : _T_53_3; // @[Mux.scala 80:57]
  wire [21:0] _T_57_3 = _T_181 ? tagArrayWire_27_3 : _T_55_3; // @[Mux.scala 80:57]
  wire [21:0] _T_59_3 = _T_183 ? tagArrayWire_28_3 : _T_57_3; // @[Mux.scala 80:57]
  wire [21:0] _T_61_3 = _T_185 ? tagArrayWire_29_3 : _T_59_3; // @[Mux.scala 80:57]
  wire [21:0] _T_63_3 = _T_187 ? tagArrayWire_30_3 : _T_61_3; // @[Mux.scala 80:57]
  wire [21:0] _T_65_3 = _T_189 ? tagArrayWire_31_3 : _T_63_3; // @[Mux.scala 80:57]
  wire [21:0] _T_67_3 = _T_191 ? tagArrayWire_32_3 : _T_65_3; // @[Mux.scala 80:57]
  wire [21:0] _T_69_3 = _T_193 ? tagArrayWire_33_3 : _T_67_3; // @[Mux.scala 80:57]
  wire [21:0] _T_71_3 = _T_195 ? tagArrayWire_34_3 : _T_69_3; // @[Mux.scala 80:57]
  wire [21:0] _T_73_3 = _T_197 ? tagArrayWire_35_3 : _T_71_3; // @[Mux.scala 80:57]
  wire [21:0] _T_75_3 = _T_199 ? tagArrayWire_36_3 : _T_73_3; // @[Mux.scala 80:57]
  wire [21:0] _T_77_3 = _T_201 ? tagArrayWire_37_3 : _T_75_3; // @[Mux.scala 80:57]
  wire [21:0] _T_79_3 = _T_203 ? tagArrayWire_38_3 : _T_77_3; // @[Mux.scala 80:57]
  wire [21:0] _T_81_3 = _T_205 ? tagArrayWire_39_3 : _T_79_3; // @[Mux.scala 80:57]
  wire [21:0] _T_83_3 = _T_207 ? tagArrayWire_40_3 : _T_81_3; // @[Mux.scala 80:57]
  wire [21:0] _T_85_3 = _T_209 ? tagArrayWire_41_3 : _T_83_3; // @[Mux.scala 80:57]
  wire [21:0] _T_87_3 = _T_211 ? tagArrayWire_42_3 : _T_85_3; // @[Mux.scala 80:57]
  wire [21:0] _T_89_3 = _T_213 ? tagArrayWire_43_3 : _T_87_3; // @[Mux.scala 80:57]
  wire [21:0] _T_91_3 = _T_215 ? tagArrayWire_44_3 : _T_89_3; // @[Mux.scala 80:57]
  wire [21:0] _T_93_3 = _T_217 ? tagArrayWire_45_3 : _T_91_3; // @[Mux.scala 80:57]
  wire [21:0] _T_95_3 = _T_219 ? tagArrayWire_46_3 : _T_93_3; // @[Mux.scala 80:57]
  wire [21:0] _T_97_3 = _T_221 ? tagArrayWire_47_3 : _T_95_3; // @[Mux.scala 80:57]
  wire [21:0] _T_99_3 = _T_223 ? tagArrayWire_48_3 : _T_97_3; // @[Mux.scala 80:57]
  wire [21:0] _T_101_3 = _T_225 ? tagArrayWire_49_3 : _T_99_3; // @[Mux.scala 80:57]
  wire [21:0] _T_103_3 = _T_227 ? tagArrayWire_50_3 : _T_101_3; // @[Mux.scala 80:57]
  wire [21:0] _T_105_3 = _T_229 ? tagArrayWire_51_3 : _T_103_3; // @[Mux.scala 80:57]
  wire [21:0] _T_107_3 = _T_231 ? tagArrayWire_52_3 : _T_105_3; // @[Mux.scala 80:57]
  wire [21:0] _T_109_3 = _T_233 ? tagArrayWire_53_3 : _T_107_3; // @[Mux.scala 80:57]
  wire [21:0] _T_111_3 = _T_235 ? tagArrayWire_54_3 : _T_109_3; // @[Mux.scala 80:57]
  wire [21:0] _T_113_3 = _T_237 ? tagArrayWire_55_3 : _T_111_3; // @[Mux.scala 80:57]
  wire [21:0] _T_115_3 = _T_239 ? tagArrayWire_56_3 : _T_113_3; // @[Mux.scala 80:57]
  wire [21:0] _T_117_3 = _T_241 ? tagArrayWire_57_3 : _T_115_3; // @[Mux.scala 80:57]
  wire [21:0] _T_119_3 = _T_243 ? tagArrayWire_58_3 : _T_117_3; // @[Mux.scala 80:57]
  wire [21:0] _T_121_3 = _T_245 ? tagArrayWire_59_3 : _T_119_3; // @[Mux.scala 80:57]
  wire [21:0] _T_123_3 = _T_247 ? tagArrayWire_60_3 : _T_121_3; // @[Mux.scala 80:57]
  wire [21:0] _T_125_3 = _T_249 ? tagArrayWire_61_3 : _T_123_3; // @[Mux.scala 80:57]
  wire [21:0] _T_127_3 = _T_251 ? tagArrayWire_62_3 : _T_125_3; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_3 = _T_253 ? tagArrayWire_63_3 : _T_127_3; // @[Mux.scala 80:57]
  wire  _T_257 = tagMuxOut_3 == tag; // @[Cache.scala 72:76]
  wire  hitArray_3 = vMuxOut_3 & _T_257; // @[Cache.scala 72:60]
  wire  hit = _T_260 | hitArray_3; // @[Cache.scala 73:49]
  wire  _T = ~hit; // @[Cache.scala 35:41]
  wire  IdleMux = io_cacheIn_valid & _T; // @[Cache.scala 35:38]
  wire  isIdle = ~cacheState; // @[Cache.scala 45:27]
  wire [127:0] _T_262 = hitArray_0 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_263 = hitArray_1 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_264 = hitArray_2 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_265 = hitArray_3 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_266 = _T_262 | _T_263; // @[Mux.scala 27:72]
  wire [127:0] _T_267 = _T_266 | _T_264; // @[Mux.scala 27:72]
  wire [127:0] waysel = _T_267 | _T_265; // @[Mux.scala 27:72]
  reg [1:0] selArrayWire_1; // @[Reg.scala 27:20]
  reg [1:0] selArrayWire_0; // @[Reg.scala 27:20]
  wire [1:0] _T_274 = _T_129 ? selArrayWire_1 : selArrayWire_0; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_2; // @[Reg.scala 27:20]
  wire [1:0] _T_276 = _T_131 ? selArrayWire_2 : _T_274; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_3; // @[Reg.scala 27:20]
  wire [1:0] _T_278 = _T_133 ? selArrayWire_3 : _T_276; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_4; // @[Reg.scala 27:20]
  wire [1:0] _T_280 = _T_135 ? selArrayWire_4 : _T_278; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_5; // @[Reg.scala 27:20]
  wire [1:0] _T_282 = _T_137 ? selArrayWire_5 : _T_280; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_6; // @[Reg.scala 27:20]
  wire [1:0] _T_284 = _T_139 ? selArrayWire_6 : _T_282; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_7; // @[Reg.scala 27:20]
  wire [1:0] _T_286 = _T_141 ? selArrayWire_7 : _T_284; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_8; // @[Reg.scala 27:20]
  wire [1:0] _T_288 = _T_143 ? selArrayWire_8 : _T_286; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_9; // @[Reg.scala 27:20]
  wire [1:0] _T_290 = _T_145 ? selArrayWire_9 : _T_288; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_10; // @[Reg.scala 27:20]
  wire [1:0] _T_292 = _T_147 ? selArrayWire_10 : _T_290; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_11; // @[Reg.scala 27:20]
  wire [1:0] _T_294 = _T_149 ? selArrayWire_11 : _T_292; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_12; // @[Reg.scala 27:20]
  wire [1:0] _T_296 = _T_151 ? selArrayWire_12 : _T_294; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_13; // @[Reg.scala 27:20]
  wire [1:0] _T_298 = _T_153 ? selArrayWire_13 : _T_296; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_14; // @[Reg.scala 27:20]
  wire [1:0] _T_300 = _T_155 ? selArrayWire_14 : _T_298; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_15; // @[Reg.scala 27:20]
  wire [1:0] _T_302 = _T_157 ? selArrayWire_15 : _T_300; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_16; // @[Reg.scala 27:20]
  wire [1:0] _T_304 = _T_159 ? selArrayWire_16 : _T_302; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_17; // @[Reg.scala 27:20]
  wire [1:0] _T_306 = _T_161 ? selArrayWire_17 : _T_304; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_18; // @[Reg.scala 27:20]
  wire [1:0] _T_308 = _T_163 ? selArrayWire_18 : _T_306; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_19; // @[Reg.scala 27:20]
  wire [1:0] _T_310 = _T_165 ? selArrayWire_19 : _T_308; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_20; // @[Reg.scala 27:20]
  wire [1:0] _T_312 = _T_167 ? selArrayWire_20 : _T_310; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_21; // @[Reg.scala 27:20]
  wire [1:0] _T_314 = _T_169 ? selArrayWire_21 : _T_312; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_22; // @[Reg.scala 27:20]
  wire [1:0] _T_316 = _T_171 ? selArrayWire_22 : _T_314; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_23; // @[Reg.scala 27:20]
  wire [1:0] _T_318 = _T_173 ? selArrayWire_23 : _T_316; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_24; // @[Reg.scala 27:20]
  wire [1:0] _T_320 = _T_175 ? selArrayWire_24 : _T_318; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_25; // @[Reg.scala 27:20]
  wire [1:0] _T_322 = _T_177 ? selArrayWire_25 : _T_320; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_26; // @[Reg.scala 27:20]
  wire [1:0] _T_324 = _T_179 ? selArrayWire_26 : _T_322; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_27; // @[Reg.scala 27:20]
  wire [1:0] _T_326 = _T_181 ? selArrayWire_27 : _T_324; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_28; // @[Reg.scala 27:20]
  wire [1:0] _T_328 = _T_183 ? selArrayWire_28 : _T_326; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_29; // @[Reg.scala 27:20]
  wire [1:0] _T_330 = _T_185 ? selArrayWire_29 : _T_328; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_30; // @[Reg.scala 27:20]
  wire [1:0] _T_332 = _T_187 ? selArrayWire_30 : _T_330; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_31; // @[Reg.scala 27:20]
  wire [1:0] _T_334 = _T_189 ? selArrayWire_31 : _T_332; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_32; // @[Reg.scala 27:20]
  wire [1:0] _T_336 = _T_191 ? selArrayWire_32 : _T_334; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_33; // @[Reg.scala 27:20]
  wire [1:0] _T_338 = _T_193 ? selArrayWire_33 : _T_336; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_34; // @[Reg.scala 27:20]
  wire [1:0] _T_340 = _T_195 ? selArrayWire_34 : _T_338; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_35; // @[Reg.scala 27:20]
  wire [1:0] _T_342 = _T_197 ? selArrayWire_35 : _T_340; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_36; // @[Reg.scala 27:20]
  wire [1:0] _T_344 = _T_199 ? selArrayWire_36 : _T_342; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_37; // @[Reg.scala 27:20]
  wire [1:0] _T_346 = _T_201 ? selArrayWire_37 : _T_344; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_38; // @[Reg.scala 27:20]
  wire [1:0] _T_348 = _T_203 ? selArrayWire_38 : _T_346; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_39; // @[Reg.scala 27:20]
  wire [1:0] _T_350 = _T_205 ? selArrayWire_39 : _T_348; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_40; // @[Reg.scala 27:20]
  wire [1:0] _T_352 = _T_207 ? selArrayWire_40 : _T_350; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_41; // @[Reg.scala 27:20]
  wire [1:0] _T_354 = _T_209 ? selArrayWire_41 : _T_352; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_42; // @[Reg.scala 27:20]
  wire [1:0] _T_356 = _T_211 ? selArrayWire_42 : _T_354; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_43; // @[Reg.scala 27:20]
  wire [1:0] _T_358 = _T_213 ? selArrayWire_43 : _T_356; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_44; // @[Reg.scala 27:20]
  wire [1:0] _T_360 = _T_215 ? selArrayWire_44 : _T_358; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_45; // @[Reg.scala 27:20]
  wire [1:0] _T_362 = _T_217 ? selArrayWire_45 : _T_360; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_46; // @[Reg.scala 27:20]
  wire [1:0] _T_364 = _T_219 ? selArrayWire_46 : _T_362; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_47; // @[Reg.scala 27:20]
  wire [1:0] _T_366 = _T_221 ? selArrayWire_47 : _T_364; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_48; // @[Reg.scala 27:20]
  wire [1:0] _T_368 = _T_223 ? selArrayWire_48 : _T_366; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_49; // @[Reg.scala 27:20]
  wire [1:0] _T_370 = _T_225 ? selArrayWire_49 : _T_368; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_50; // @[Reg.scala 27:20]
  wire [1:0] _T_372 = _T_227 ? selArrayWire_50 : _T_370; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_51; // @[Reg.scala 27:20]
  wire [1:0] _T_374 = _T_229 ? selArrayWire_51 : _T_372; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_52; // @[Reg.scala 27:20]
  wire [1:0] _T_376 = _T_231 ? selArrayWire_52 : _T_374; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_53; // @[Reg.scala 27:20]
  wire [1:0] _T_378 = _T_233 ? selArrayWire_53 : _T_376; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_54; // @[Reg.scala 27:20]
  wire [1:0] _T_380 = _T_235 ? selArrayWire_54 : _T_378; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_55; // @[Reg.scala 27:20]
  wire [1:0] _T_382 = _T_237 ? selArrayWire_55 : _T_380; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_56; // @[Reg.scala 27:20]
  wire [1:0] _T_384 = _T_239 ? selArrayWire_56 : _T_382; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_57; // @[Reg.scala 27:20]
  wire [1:0] _T_386 = _T_241 ? selArrayWire_57 : _T_384; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_58; // @[Reg.scala 27:20]
  wire [1:0] _T_388 = _T_243 ? selArrayWire_58 : _T_386; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_59; // @[Reg.scala 27:20]
  wire [1:0] _T_390 = _T_245 ? selArrayWire_59 : _T_388; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_60; // @[Reg.scala 27:20]
  wire [1:0] _T_392 = _T_247 ? selArrayWire_60 : _T_390; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_61; // @[Reg.scala 27:20]
  wire [1:0] _T_394 = _T_249 ? selArrayWire_61 : _T_392; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_62; // @[Reg.scala 27:20]
  wire [1:0] _T_396 = _T_251 ? selArrayWire_62 : _T_394; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_63; // @[Reg.scala 27:20]
  wire [1:0] sramSel = _T_253 ? selArrayWire_63 : _T_396; // @[Mux.scala 80:57]
  wire [1:0] _T_401 = selArrayWire_0 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_402 = 6'h0 == index; // @[Cache.scala 111:36]
  wire  _T_403 = io_cacheOut_r_last_i & _T_402; // @[Cache.scala 111:28]
  wire  _T_407 = selArrayWire_0 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_408 = _T_403 & _T_407; // @[Cache.scala 114:85]
  wire  _T_409 = _T_408 & cacheState; // @[Cache.scala 114:112]
  wire  _T_412 = reset | updataICache_0; // @[Cache.scala 115:33]
  wire  _GEN_2 = _T_409 | vArrayWire_0_0; // @[Reg.scala 28:19]
  wire  _T_421 = selArrayWire_0 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_422 = _T_403 & _T_421; // @[Cache.scala 114:85]
  wire  _T_423 = _T_422 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_4 = _T_423 | vArrayWire_0_1; // @[Reg.scala 28:19]
  wire  _T_435 = selArrayWire_0 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_436 = _T_403 & _T_435; // @[Cache.scala 114:85]
  wire  _T_437 = _T_436 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_6 = _T_437 | vArrayWire_0_2; // @[Reg.scala 28:19]
  wire  _T_449 = selArrayWire_0 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_450 = _T_403 & _T_449; // @[Cache.scala 114:85]
  wire  _T_451 = _T_450 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_8 = _T_451 | vArrayWire_0_3; // @[Reg.scala 28:19]
  wire [1:0] _T_462 = selArrayWire_1 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_464 = io_cacheOut_r_last_i & _T_129; // @[Cache.scala 111:28]
  wire  _T_468 = selArrayWire_1 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_469 = _T_464 & _T_468; // @[Cache.scala 114:85]
  wire  _T_470 = _T_469 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_11 = _T_470 | vArrayWire_1_0; // @[Reg.scala 28:19]
  wire  _T_482 = selArrayWire_1 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_483 = _T_464 & _T_482; // @[Cache.scala 114:85]
  wire  _T_484 = _T_483 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_13 = _T_484 | vArrayWire_1_1; // @[Reg.scala 28:19]
  wire  _T_496 = selArrayWire_1 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_497 = _T_464 & _T_496; // @[Cache.scala 114:85]
  wire  _T_498 = _T_497 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_15 = _T_498 | vArrayWire_1_2; // @[Reg.scala 28:19]
  wire  _T_510 = selArrayWire_1 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_511 = _T_464 & _T_510; // @[Cache.scala 114:85]
  wire  _T_512 = _T_511 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_17 = _T_512 | vArrayWire_1_3; // @[Reg.scala 28:19]
  wire [1:0] _T_523 = selArrayWire_2 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_525 = io_cacheOut_r_last_i & _T_131; // @[Cache.scala 111:28]
  wire  _T_529 = selArrayWire_2 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_530 = _T_525 & _T_529; // @[Cache.scala 114:85]
  wire  _T_531 = _T_530 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_20 = _T_531 | vArrayWire_2_0; // @[Reg.scala 28:19]
  wire  _T_543 = selArrayWire_2 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_544 = _T_525 & _T_543; // @[Cache.scala 114:85]
  wire  _T_545 = _T_544 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_22 = _T_545 | vArrayWire_2_1; // @[Reg.scala 28:19]
  wire  _T_557 = selArrayWire_2 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_558 = _T_525 & _T_557; // @[Cache.scala 114:85]
  wire  _T_559 = _T_558 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_24 = _T_559 | vArrayWire_2_2; // @[Reg.scala 28:19]
  wire  _T_571 = selArrayWire_2 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_572 = _T_525 & _T_571; // @[Cache.scala 114:85]
  wire  _T_573 = _T_572 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_26 = _T_573 | vArrayWire_2_3; // @[Reg.scala 28:19]
  wire [1:0] _T_584 = selArrayWire_3 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_586 = io_cacheOut_r_last_i & _T_133; // @[Cache.scala 111:28]
  wire  _T_590 = selArrayWire_3 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_591 = _T_586 & _T_590; // @[Cache.scala 114:85]
  wire  _T_592 = _T_591 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_29 = _T_592 | vArrayWire_3_0; // @[Reg.scala 28:19]
  wire  _T_604 = selArrayWire_3 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_605 = _T_586 & _T_604; // @[Cache.scala 114:85]
  wire  _T_606 = _T_605 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_31 = _T_606 | vArrayWire_3_1; // @[Reg.scala 28:19]
  wire  _T_618 = selArrayWire_3 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_619 = _T_586 & _T_618; // @[Cache.scala 114:85]
  wire  _T_620 = _T_619 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_33 = _T_620 | vArrayWire_3_2; // @[Reg.scala 28:19]
  wire  _T_632 = selArrayWire_3 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_633 = _T_586 & _T_632; // @[Cache.scala 114:85]
  wire  _T_634 = _T_633 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_35 = _T_634 | vArrayWire_3_3; // @[Reg.scala 28:19]
  wire [1:0] _T_645 = selArrayWire_4 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_647 = io_cacheOut_r_last_i & _T_135; // @[Cache.scala 111:28]
  wire  _T_651 = selArrayWire_4 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_652 = _T_647 & _T_651; // @[Cache.scala 114:85]
  wire  _T_653 = _T_652 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_38 = _T_653 | vArrayWire_4_0; // @[Reg.scala 28:19]
  wire  _T_665 = selArrayWire_4 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_666 = _T_647 & _T_665; // @[Cache.scala 114:85]
  wire  _T_667 = _T_666 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_40 = _T_667 | vArrayWire_4_1; // @[Reg.scala 28:19]
  wire  _T_679 = selArrayWire_4 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_680 = _T_647 & _T_679; // @[Cache.scala 114:85]
  wire  _T_681 = _T_680 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_42 = _T_681 | vArrayWire_4_2; // @[Reg.scala 28:19]
  wire  _T_693 = selArrayWire_4 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_694 = _T_647 & _T_693; // @[Cache.scala 114:85]
  wire  _T_695 = _T_694 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_44 = _T_695 | vArrayWire_4_3; // @[Reg.scala 28:19]
  wire [1:0] _T_706 = selArrayWire_5 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_708 = io_cacheOut_r_last_i & _T_137; // @[Cache.scala 111:28]
  wire  _T_712 = selArrayWire_5 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_713 = _T_708 & _T_712; // @[Cache.scala 114:85]
  wire  _T_714 = _T_713 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_47 = _T_714 | vArrayWire_5_0; // @[Reg.scala 28:19]
  wire  _T_726 = selArrayWire_5 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_727 = _T_708 & _T_726; // @[Cache.scala 114:85]
  wire  _T_728 = _T_727 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_49 = _T_728 | vArrayWire_5_1; // @[Reg.scala 28:19]
  wire  _T_740 = selArrayWire_5 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_741 = _T_708 & _T_740; // @[Cache.scala 114:85]
  wire  _T_742 = _T_741 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_51 = _T_742 | vArrayWire_5_2; // @[Reg.scala 28:19]
  wire  _T_754 = selArrayWire_5 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_755 = _T_708 & _T_754; // @[Cache.scala 114:85]
  wire  _T_756 = _T_755 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_53 = _T_756 | vArrayWire_5_3; // @[Reg.scala 28:19]
  wire [1:0] _T_767 = selArrayWire_6 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_769 = io_cacheOut_r_last_i & _T_139; // @[Cache.scala 111:28]
  wire  _T_773 = selArrayWire_6 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_774 = _T_769 & _T_773; // @[Cache.scala 114:85]
  wire  _T_775 = _T_774 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_56 = _T_775 | vArrayWire_6_0; // @[Reg.scala 28:19]
  wire  _T_787 = selArrayWire_6 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_788 = _T_769 & _T_787; // @[Cache.scala 114:85]
  wire  _T_789 = _T_788 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_58 = _T_789 | vArrayWire_6_1; // @[Reg.scala 28:19]
  wire  _T_801 = selArrayWire_6 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_802 = _T_769 & _T_801; // @[Cache.scala 114:85]
  wire  _T_803 = _T_802 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_60 = _T_803 | vArrayWire_6_2; // @[Reg.scala 28:19]
  wire  _T_815 = selArrayWire_6 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_816 = _T_769 & _T_815; // @[Cache.scala 114:85]
  wire  _T_817 = _T_816 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_62 = _T_817 | vArrayWire_6_3; // @[Reg.scala 28:19]
  wire [1:0] _T_828 = selArrayWire_7 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_830 = io_cacheOut_r_last_i & _T_141; // @[Cache.scala 111:28]
  wire  _T_834 = selArrayWire_7 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_835 = _T_830 & _T_834; // @[Cache.scala 114:85]
  wire  _T_836 = _T_835 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_65 = _T_836 | vArrayWire_7_0; // @[Reg.scala 28:19]
  wire  _T_848 = selArrayWire_7 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_849 = _T_830 & _T_848; // @[Cache.scala 114:85]
  wire  _T_850 = _T_849 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_67 = _T_850 | vArrayWire_7_1; // @[Reg.scala 28:19]
  wire  _T_862 = selArrayWire_7 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_863 = _T_830 & _T_862; // @[Cache.scala 114:85]
  wire  _T_864 = _T_863 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_69 = _T_864 | vArrayWire_7_2; // @[Reg.scala 28:19]
  wire  _T_876 = selArrayWire_7 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_877 = _T_830 & _T_876; // @[Cache.scala 114:85]
  wire  _T_878 = _T_877 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_71 = _T_878 | vArrayWire_7_3; // @[Reg.scala 28:19]
  wire [1:0] _T_889 = selArrayWire_8 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_891 = io_cacheOut_r_last_i & _T_143; // @[Cache.scala 111:28]
  wire  _T_895 = selArrayWire_8 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_896 = _T_891 & _T_895; // @[Cache.scala 114:85]
  wire  _T_897 = _T_896 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_74 = _T_897 | vArrayWire_8_0; // @[Reg.scala 28:19]
  wire  _T_909 = selArrayWire_8 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_910 = _T_891 & _T_909; // @[Cache.scala 114:85]
  wire  _T_911 = _T_910 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_76 = _T_911 | vArrayWire_8_1; // @[Reg.scala 28:19]
  wire  _T_923 = selArrayWire_8 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_924 = _T_891 & _T_923; // @[Cache.scala 114:85]
  wire  _T_925 = _T_924 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_78 = _T_925 | vArrayWire_8_2; // @[Reg.scala 28:19]
  wire  _T_937 = selArrayWire_8 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_938 = _T_891 & _T_937; // @[Cache.scala 114:85]
  wire  _T_939 = _T_938 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_80 = _T_939 | vArrayWire_8_3; // @[Reg.scala 28:19]
  wire [1:0] _T_950 = selArrayWire_9 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_952 = io_cacheOut_r_last_i & _T_145; // @[Cache.scala 111:28]
  wire  _T_956 = selArrayWire_9 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_957 = _T_952 & _T_956; // @[Cache.scala 114:85]
  wire  _T_958 = _T_957 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_83 = _T_958 | vArrayWire_9_0; // @[Reg.scala 28:19]
  wire  _T_970 = selArrayWire_9 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_971 = _T_952 & _T_970; // @[Cache.scala 114:85]
  wire  _T_972 = _T_971 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_85 = _T_972 | vArrayWire_9_1; // @[Reg.scala 28:19]
  wire  _T_984 = selArrayWire_9 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_985 = _T_952 & _T_984; // @[Cache.scala 114:85]
  wire  _T_986 = _T_985 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_87 = _T_986 | vArrayWire_9_2; // @[Reg.scala 28:19]
  wire  _T_998 = selArrayWire_9 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_999 = _T_952 & _T_998; // @[Cache.scala 114:85]
  wire  _T_1000 = _T_999 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_89 = _T_1000 | vArrayWire_9_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1011 = selArrayWire_10 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1013 = io_cacheOut_r_last_i & _T_147; // @[Cache.scala 111:28]
  wire  _T_1017 = selArrayWire_10 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1018 = _T_1013 & _T_1017; // @[Cache.scala 114:85]
  wire  _T_1019 = _T_1018 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_92 = _T_1019 | vArrayWire_10_0; // @[Reg.scala 28:19]
  wire  _T_1031 = selArrayWire_10 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1032 = _T_1013 & _T_1031; // @[Cache.scala 114:85]
  wire  _T_1033 = _T_1032 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_94 = _T_1033 | vArrayWire_10_1; // @[Reg.scala 28:19]
  wire  _T_1045 = selArrayWire_10 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1046 = _T_1013 & _T_1045; // @[Cache.scala 114:85]
  wire  _T_1047 = _T_1046 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_96 = _T_1047 | vArrayWire_10_2; // @[Reg.scala 28:19]
  wire  _T_1059 = selArrayWire_10 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1060 = _T_1013 & _T_1059; // @[Cache.scala 114:85]
  wire  _T_1061 = _T_1060 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_98 = _T_1061 | vArrayWire_10_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1072 = selArrayWire_11 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1074 = io_cacheOut_r_last_i & _T_149; // @[Cache.scala 111:28]
  wire  _T_1078 = selArrayWire_11 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1079 = _T_1074 & _T_1078; // @[Cache.scala 114:85]
  wire  _T_1080 = _T_1079 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_101 = _T_1080 | vArrayWire_11_0; // @[Reg.scala 28:19]
  wire  _T_1092 = selArrayWire_11 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1093 = _T_1074 & _T_1092; // @[Cache.scala 114:85]
  wire  _T_1094 = _T_1093 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_103 = _T_1094 | vArrayWire_11_1; // @[Reg.scala 28:19]
  wire  _T_1106 = selArrayWire_11 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1107 = _T_1074 & _T_1106; // @[Cache.scala 114:85]
  wire  _T_1108 = _T_1107 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_105 = _T_1108 | vArrayWire_11_2; // @[Reg.scala 28:19]
  wire  _T_1120 = selArrayWire_11 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1121 = _T_1074 & _T_1120; // @[Cache.scala 114:85]
  wire  _T_1122 = _T_1121 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_107 = _T_1122 | vArrayWire_11_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1133 = selArrayWire_12 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1135 = io_cacheOut_r_last_i & _T_151; // @[Cache.scala 111:28]
  wire  _T_1139 = selArrayWire_12 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1140 = _T_1135 & _T_1139; // @[Cache.scala 114:85]
  wire  _T_1141 = _T_1140 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_110 = _T_1141 | vArrayWire_12_0; // @[Reg.scala 28:19]
  wire  _T_1153 = selArrayWire_12 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1154 = _T_1135 & _T_1153; // @[Cache.scala 114:85]
  wire  _T_1155 = _T_1154 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_112 = _T_1155 | vArrayWire_12_1; // @[Reg.scala 28:19]
  wire  _T_1167 = selArrayWire_12 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1168 = _T_1135 & _T_1167; // @[Cache.scala 114:85]
  wire  _T_1169 = _T_1168 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_114 = _T_1169 | vArrayWire_12_2; // @[Reg.scala 28:19]
  wire  _T_1181 = selArrayWire_12 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1182 = _T_1135 & _T_1181; // @[Cache.scala 114:85]
  wire  _T_1183 = _T_1182 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_116 = _T_1183 | vArrayWire_12_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1194 = selArrayWire_13 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1196 = io_cacheOut_r_last_i & _T_153; // @[Cache.scala 111:28]
  wire  _T_1200 = selArrayWire_13 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1201 = _T_1196 & _T_1200; // @[Cache.scala 114:85]
  wire  _T_1202 = _T_1201 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_119 = _T_1202 | vArrayWire_13_0; // @[Reg.scala 28:19]
  wire  _T_1214 = selArrayWire_13 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1215 = _T_1196 & _T_1214; // @[Cache.scala 114:85]
  wire  _T_1216 = _T_1215 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_121 = _T_1216 | vArrayWire_13_1; // @[Reg.scala 28:19]
  wire  _T_1228 = selArrayWire_13 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1229 = _T_1196 & _T_1228; // @[Cache.scala 114:85]
  wire  _T_1230 = _T_1229 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_123 = _T_1230 | vArrayWire_13_2; // @[Reg.scala 28:19]
  wire  _T_1242 = selArrayWire_13 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1243 = _T_1196 & _T_1242; // @[Cache.scala 114:85]
  wire  _T_1244 = _T_1243 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_125 = _T_1244 | vArrayWire_13_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1255 = selArrayWire_14 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1257 = io_cacheOut_r_last_i & _T_155; // @[Cache.scala 111:28]
  wire  _T_1261 = selArrayWire_14 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1262 = _T_1257 & _T_1261; // @[Cache.scala 114:85]
  wire  _T_1263 = _T_1262 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_128 = _T_1263 | vArrayWire_14_0; // @[Reg.scala 28:19]
  wire  _T_1275 = selArrayWire_14 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1276 = _T_1257 & _T_1275; // @[Cache.scala 114:85]
  wire  _T_1277 = _T_1276 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_130 = _T_1277 | vArrayWire_14_1; // @[Reg.scala 28:19]
  wire  _T_1289 = selArrayWire_14 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1290 = _T_1257 & _T_1289; // @[Cache.scala 114:85]
  wire  _T_1291 = _T_1290 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_132 = _T_1291 | vArrayWire_14_2; // @[Reg.scala 28:19]
  wire  _T_1303 = selArrayWire_14 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1304 = _T_1257 & _T_1303; // @[Cache.scala 114:85]
  wire  _T_1305 = _T_1304 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_134 = _T_1305 | vArrayWire_14_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1316 = selArrayWire_15 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1318 = io_cacheOut_r_last_i & _T_157; // @[Cache.scala 111:28]
  wire  _T_1322 = selArrayWire_15 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1323 = _T_1318 & _T_1322; // @[Cache.scala 114:85]
  wire  _T_1324 = _T_1323 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_137 = _T_1324 | vArrayWire_15_0; // @[Reg.scala 28:19]
  wire  _T_1336 = selArrayWire_15 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1337 = _T_1318 & _T_1336; // @[Cache.scala 114:85]
  wire  _T_1338 = _T_1337 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_139 = _T_1338 | vArrayWire_15_1; // @[Reg.scala 28:19]
  wire  _T_1350 = selArrayWire_15 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1351 = _T_1318 & _T_1350; // @[Cache.scala 114:85]
  wire  _T_1352 = _T_1351 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_141 = _T_1352 | vArrayWire_15_2; // @[Reg.scala 28:19]
  wire  _T_1364 = selArrayWire_15 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1365 = _T_1318 & _T_1364; // @[Cache.scala 114:85]
  wire  _T_1366 = _T_1365 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_143 = _T_1366 | vArrayWire_15_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1377 = selArrayWire_16 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1379 = io_cacheOut_r_last_i & _T_159; // @[Cache.scala 111:28]
  wire  _T_1383 = selArrayWire_16 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1384 = _T_1379 & _T_1383; // @[Cache.scala 114:85]
  wire  _T_1385 = _T_1384 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_146 = _T_1385 | vArrayWire_16_0; // @[Reg.scala 28:19]
  wire  _T_1397 = selArrayWire_16 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1398 = _T_1379 & _T_1397; // @[Cache.scala 114:85]
  wire  _T_1399 = _T_1398 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_148 = _T_1399 | vArrayWire_16_1; // @[Reg.scala 28:19]
  wire  _T_1411 = selArrayWire_16 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1412 = _T_1379 & _T_1411; // @[Cache.scala 114:85]
  wire  _T_1413 = _T_1412 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_150 = _T_1413 | vArrayWire_16_2; // @[Reg.scala 28:19]
  wire  _T_1425 = selArrayWire_16 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1426 = _T_1379 & _T_1425; // @[Cache.scala 114:85]
  wire  _T_1427 = _T_1426 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_152 = _T_1427 | vArrayWire_16_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1438 = selArrayWire_17 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1440 = io_cacheOut_r_last_i & _T_161; // @[Cache.scala 111:28]
  wire  _T_1444 = selArrayWire_17 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1445 = _T_1440 & _T_1444; // @[Cache.scala 114:85]
  wire  _T_1446 = _T_1445 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_155 = _T_1446 | vArrayWire_17_0; // @[Reg.scala 28:19]
  wire  _T_1458 = selArrayWire_17 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1459 = _T_1440 & _T_1458; // @[Cache.scala 114:85]
  wire  _T_1460 = _T_1459 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_157 = _T_1460 | vArrayWire_17_1; // @[Reg.scala 28:19]
  wire  _T_1472 = selArrayWire_17 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1473 = _T_1440 & _T_1472; // @[Cache.scala 114:85]
  wire  _T_1474 = _T_1473 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_159 = _T_1474 | vArrayWire_17_2; // @[Reg.scala 28:19]
  wire  _T_1486 = selArrayWire_17 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1487 = _T_1440 & _T_1486; // @[Cache.scala 114:85]
  wire  _T_1488 = _T_1487 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_161 = _T_1488 | vArrayWire_17_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1499 = selArrayWire_18 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1501 = io_cacheOut_r_last_i & _T_163; // @[Cache.scala 111:28]
  wire  _T_1505 = selArrayWire_18 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1506 = _T_1501 & _T_1505; // @[Cache.scala 114:85]
  wire  _T_1507 = _T_1506 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_164 = _T_1507 | vArrayWire_18_0; // @[Reg.scala 28:19]
  wire  _T_1519 = selArrayWire_18 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1520 = _T_1501 & _T_1519; // @[Cache.scala 114:85]
  wire  _T_1521 = _T_1520 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_166 = _T_1521 | vArrayWire_18_1; // @[Reg.scala 28:19]
  wire  _T_1533 = selArrayWire_18 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1534 = _T_1501 & _T_1533; // @[Cache.scala 114:85]
  wire  _T_1535 = _T_1534 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_168 = _T_1535 | vArrayWire_18_2; // @[Reg.scala 28:19]
  wire  _T_1547 = selArrayWire_18 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1548 = _T_1501 & _T_1547; // @[Cache.scala 114:85]
  wire  _T_1549 = _T_1548 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_170 = _T_1549 | vArrayWire_18_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1560 = selArrayWire_19 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1562 = io_cacheOut_r_last_i & _T_165; // @[Cache.scala 111:28]
  wire  _T_1566 = selArrayWire_19 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1567 = _T_1562 & _T_1566; // @[Cache.scala 114:85]
  wire  _T_1568 = _T_1567 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_173 = _T_1568 | vArrayWire_19_0; // @[Reg.scala 28:19]
  wire  _T_1580 = selArrayWire_19 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1581 = _T_1562 & _T_1580; // @[Cache.scala 114:85]
  wire  _T_1582 = _T_1581 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_175 = _T_1582 | vArrayWire_19_1; // @[Reg.scala 28:19]
  wire  _T_1594 = selArrayWire_19 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1595 = _T_1562 & _T_1594; // @[Cache.scala 114:85]
  wire  _T_1596 = _T_1595 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_177 = _T_1596 | vArrayWire_19_2; // @[Reg.scala 28:19]
  wire  _T_1608 = selArrayWire_19 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1609 = _T_1562 & _T_1608; // @[Cache.scala 114:85]
  wire  _T_1610 = _T_1609 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_179 = _T_1610 | vArrayWire_19_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1621 = selArrayWire_20 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1623 = io_cacheOut_r_last_i & _T_167; // @[Cache.scala 111:28]
  wire  _T_1627 = selArrayWire_20 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1628 = _T_1623 & _T_1627; // @[Cache.scala 114:85]
  wire  _T_1629 = _T_1628 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_182 = _T_1629 | vArrayWire_20_0; // @[Reg.scala 28:19]
  wire  _T_1641 = selArrayWire_20 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1642 = _T_1623 & _T_1641; // @[Cache.scala 114:85]
  wire  _T_1643 = _T_1642 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_184 = _T_1643 | vArrayWire_20_1; // @[Reg.scala 28:19]
  wire  _T_1655 = selArrayWire_20 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1656 = _T_1623 & _T_1655; // @[Cache.scala 114:85]
  wire  _T_1657 = _T_1656 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_186 = _T_1657 | vArrayWire_20_2; // @[Reg.scala 28:19]
  wire  _T_1669 = selArrayWire_20 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1670 = _T_1623 & _T_1669; // @[Cache.scala 114:85]
  wire  _T_1671 = _T_1670 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_188 = _T_1671 | vArrayWire_20_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1682 = selArrayWire_21 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1684 = io_cacheOut_r_last_i & _T_169; // @[Cache.scala 111:28]
  wire  _T_1688 = selArrayWire_21 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1689 = _T_1684 & _T_1688; // @[Cache.scala 114:85]
  wire  _T_1690 = _T_1689 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_191 = _T_1690 | vArrayWire_21_0; // @[Reg.scala 28:19]
  wire  _T_1702 = selArrayWire_21 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1703 = _T_1684 & _T_1702; // @[Cache.scala 114:85]
  wire  _T_1704 = _T_1703 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_193 = _T_1704 | vArrayWire_21_1; // @[Reg.scala 28:19]
  wire  _T_1716 = selArrayWire_21 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1717 = _T_1684 & _T_1716; // @[Cache.scala 114:85]
  wire  _T_1718 = _T_1717 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_195 = _T_1718 | vArrayWire_21_2; // @[Reg.scala 28:19]
  wire  _T_1730 = selArrayWire_21 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1731 = _T_1684 & _T_1730; // @[Cache.scala 114:85]
  wire  _T_1732 = _T_1731 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_197 = _T_1732 | vArrayWire_21_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1743 = selArrayWire_22 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1745 = io_cacheOut_r_last_i & _T_171; // @[Cache.scala 111:28]
  wire  _T_1749 = selArrayWire_22 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1750 = _T_1745 & _T_1749; // @[Cache.scala 114:85]
  wire  _T_1751 = _T_1750 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_200 = _T_1751 | vArrayWire_22_0; // @[Reg.scala 28:19]
  wire  _T_1763 = selArrayWire_22 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1764 = _T_1745 & _T_1763; // @[Cache.scala 114:85]
  wire  _T_1765 = _T_1764 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_202 = _T_1765 | vArrayWire_22_1; // @[Reg.scala 28:19]
  wire  _T_1777 = selArrayWire_22 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1778 = _T_1745 & _T_1777; // @[Cache.scala 114:85]
  wire  _T_1779 = _T_1778 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_204 = _T_1779 | vArrayWire_22_2; // @[Reg.scala 28:19]
  wire  _T_1791 = selArrayWire_22 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1792 = _T_1745 & _T_1791; // @[Cache.scala 114:85]
  wire  _T_1793 = _T_1792 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_206 = _T_1793 | vArrayWire_22_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1804 = selArrayWire_23 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1806 = io_cacheOut_r_last_i & _T_173; // @[Cache.scala 111:28]
  wire  _T_1810 = selArrayWire_23 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1811 = _T_1806 & _T_1810; // @[Cache.scala 114:85]
  wire  _T_1812 = _T_1811 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_209 = _T_1812 | vArrayWire_23_0; // @[Reg.scala 28:19]
  wire  _T_1824 = selArrayWire_23 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1825 = _T_1806 & _T_1824; // @[Cache.scala 114:85]
  wire  _T_1826 = _T_1825 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_211 = _T_1826 | vArrayWire_23_1; // @[Reg.scala 28:19]
  wire  _T_1838 = selArrayWire_23 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1839 = _T_1806 & _T_1838; // @[Cache.scala 114:85]
  wire  _T_1840 = _T_1839 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_213 = _T_1840 | vArrayWire_23_2; // @[Reg.scala 28:19]
  wire  _T_1852 = selArrayWire_23 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1853 = _T_1806 & _T_1852; // @[Cache.scala 114:85]
  wire  _T_1854 = _T_1853 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_215 = _T_1854 | vArrayWire_23_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1865 = selArrayWire_24 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1867 = io_cacheOut_r_last_i & _T_175; // @[Cache.scala 111:28]
  wire  _T_1871 = selArrayWire_24 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1872 = _T_1867 & _T_1871; // @[Cache.scala 114:85]
  wire  _T_1873 = _T_1872 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_218 = _T_1873 | vArrayWire_24_0; // @[Reg.scala 28:19]
  wire  _T_1885 = selArrayWire_24 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1886 = _T_1867 & _T_1885; // @[Cache.scala 114:85]
  wire  _T_1887 = _T_1886 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_220 = _T_1887 | vArrayWire_24_1; // @[Reg.scala 28:19]
  wire  _T_1899 = selArrayWire_24 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1900 = _T_1867 & _T_1899; // @[Cache.scala 114:85]
  wire  _T_1901 = _T_1900 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_222 = _T_1901 | vArrayWire_24_2; // @[Reg.scala 28:19]
  wire  _T_1913 = selArrayWire_24 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1914 = _T_1867 & _T_1913; // @[Cache.scala 114:85]
  wire  _T_1915 = _T_1914 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_224 = _T_1915 | vArrayWire_24_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1926 = selArrayWire_25 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1928 = io_cacheOut_r_last_i & _T_177; // @[Cache.scala 111:28]
  wire  _T_1932 = selArrayWire_25 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1933 = _T_1928 & _T_1932; // @[Cache.scala 114:85]
  wire  _T_1934 = _T_1933 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_227 = _T_1934 | vArrayWire_25_0; // @[Reg.scala 28:19]
  wire  _T_1946 = selArrayWire_25 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_1947 = _T_1928 & _T_1946; // @[Cache.scala 114:85]
  wire  _T_1948 = _T_1947 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_229 = _T_1948 | vArrayWire_25_1; // @[Reg.scala 28:19]
  wire  _T_1960 = selArrayWire_25 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_1961 = _T_1928 & _T_1960; // @[Cache.scala 114:85]
  wire  _T_1962 = _T_1961 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_231 = _T_1962 | vArrayWire_25_2; // @[Reg.scala 28:19]
  wire  _T_1974 = selArrayWire_25 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_1975 = _T_1928 & _T_1974; // @[Cache.scala 114:85]
  wire  _T_1976 = _T_1975 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_233 = _T_1976 | vArrayWire_25_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1987 = selArrayWire_26 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_1989 = io_cacheOut_r_last_i & _T_179; // @[Cache.scala 111:28]
  wire  _T_1993 = selArrayWire_26 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_1994 = _T_1989 & _T_1993; // @[Cache.scala 114:85]
  wire  _T_1995 = _T_1994 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_236 = _T_1995 | vArrayWire_26_0; // @[Reg.scala 28:19]
  wire  _T_2007 = selArrayWire_26 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2008 = _T_1989 & _T_2007; // @[Cache.scala 114:85]
  wire  _T_2009 = _T_2008 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_238 = _T_2009 | vArrayWire_26_1; // @[Reg.scala 28:19]
  wire  _T_2021 = selArrayWire_26 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2022 = _T_1989 & _T_2021; // @[Cache.scala 114:85]
  wire  _T_2023 = _T_2022 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_240 = _T_2023 | vArrayWire_26_2; // @[Reg.scala 28:19]
  wire  _T_2035 = selArrayWire_26 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2036 = _T_1989 & _T_2035; // @[Cache.scala 114:85]
  wire  _T_2037 = _T_2036 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_242 = _T_2037 | vArrayWire_26_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2048 = selArrayWire_27 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2050 = io_cacheOut_r_last_i & _T_181; // @[Cache.scala 111:28]
  wire  _T_2054 = selArrayWire_27 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2055 = _T_2050 & _T_2054; // @[Cache.scala 114:85]
  wire  _T_2056 = _T_2055 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_245 = _T_2056 | vArrayWire_27_0; // @[Reg.scala 28:19]
  wire  _T_2068 = selArrayWire_27 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2069 = _T_2050 & _T_2068; // @[Cache.scala 114:85]
  wire  _T_2070 = _T_2069 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_247 = _T_2070 | vArrayWire_27_1; // @[Reg.scala 28:19]
  wire  _T_2082 = selArrayWire_27 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2083 = _T_2050 & _T_2082; // @[Cache.scala 114:85]
  wire  _T_2084 = _T_2083 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_249 = _T_2084 | vArrayWire_27_2; // @[Reg.scala 28:19]
  wire  _T_2096 = selArrayWire_27 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2097 = _T_2050 & _T_2096; // @[Cache.scala 114:85]
  wire  _T_2098 = _T_2097 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_251 = _T_2098 | vArrayWire_27_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2109 = selArrayWire_28 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2111 = io_cacheOut_r_last_i & _T_183; // @[Cache.scala 111:28]
  wire  _T_2115 = selArrayWire_28 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2116 = _T_2111 & _T_2115; // @[Cache.scala 114:85]
  wire  _T_2117 = _T_2116 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_254 = _T_2117 | vArrayWire_28_0; // @[Reg.scala 28:19]
  wire  _T_2129 = selArrayWire_28 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2130 = _T_2111 & _T_2129; // @[Cache.scala 114:85]
  wire  _T_2131 = _T_2130 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_256 = _T_2131 | vArrayWire_28_1; // @[Reg.scala 28:19]
  wire  _T_2143 = selArrayWire_28 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2144 = _T_2111 & _T_2143; // @[Cache.scala 114:85]
  wire  _T_2145 = _T_2144 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_258 = _T_2145 | vArrayWire_28_2; // @[Reg.scala 28:19]
  wire  _T_2157 = selArrayWire_28 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2158 = _T_2111 & _T_2157; // @[Cache.scala 114:85]
  wire  _T_2159 = _T_2158 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_260 = _T_2159 | vArrayWire_28_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2170 = selArrayWire_29 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2172 = io_cacheOut_r_last_i & _T_185; // @[Cache.scala 111:28]
  wire  _T_2176 = selArrayWire_29 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2177 = _T_2172 & _T_2176; // @[Cache.scala 114:85]
  wire  _T_2178 = _T_2177 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_263 = _T_2178 | vArrayWire_29_0; // @[Reg.scala 28:19]
  wire  _T_2190 = selArrayWire_29 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2191 = _T_2172 & _T_2190; // @[Cache.scala 114:85]
  wire  _T_2192 = _T_2191 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_265 = _T_2192 | vArrayWire_29_1; // @[Reg.scala 28:19]
  wire  _T_2204 = selArrayWire_29 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2205 = _T_2172 & _T_2204; // @[Cache.scala 114:85]
  wire  _T_2206 = _T_2205 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_267 = _T_2206 | vArrayWire_29_2; // @[Reg.scala 28:19]
  wire  _T_2218 = selArrayWire_29 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2219 = _T_2172 & _T_2218; // @[Cache.scala 114:85]
  wire  _T_2220 = _T_2219 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_269 = _T_2220 | vArrayWire_29_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2231 = selArrayWire_30 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2233 = io_cacheOut_r_last_i & _T_187; // @[Cache.scala 111:28]
  wire  _T_2237 = selArrayWire_30 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2238 = _T_2233 & _T_2237; // @[Cache.scala 114:85]
  wire  _T_2239 = _T_2238 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_272 = _T_2239 | vArrayWire_30_0; // @[Reg.scala 28:19]
  wire  _T_2251 = selArrayWire_30 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2252 = _T_2233 & _T_2251; // @[Cache.scala 114:85]
  wire  _T_2253 = _T_2252 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_274 = _T_2253 | vArrayWire_30_1; // @[Reg.scala 28:19]
  wire  _T_2265 = selArrayWire_30 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2266 = _T_2233 & _T_2265; // @[Cache.scala 114:85]
  wire  _T_2267 = _T_2266 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_276 = _T_2267 | vArrayWire_30_2; // @[Reg.scala 28:19]
  wire  _T_2279 = selArrayWire_30 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2280 = _T_2233 & _T_2279; // @[Cache.scala 114:85]
  wire  _T_2281 = _T_2280 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_278 = _T_2281 | vArrayWire_30_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2292 = selArrayWire_31 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2294 = io_cacheOut_r_last_i & _T_189; // @[Cache.scala 111:28]
  wire  _T_2298 = selArrayWire_31 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2299 = _T_2294 & _T_2298; // @[Cache.scala 114:85]
  wire  _T_2300 = _T_2299 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_281 = _T_2300 | vArrayWire_31_0; // @[Reg.scala 28:19]
  wire  _T_2312 = selArrayWire_31 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2313 = _T_2294 & _T_2312; // @[Cache.scala 114:85]
  wire  _T_2314 = _T_2313 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_283 = _T_2314 | vArrayWire_31_1; // @[Reg.scala 28:19]
  wire  _T_2326 = selArrayWire_31 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2327 = _T_2294 & _T_2326; // @[Cache.scala 114:85]
  wire  _T_2328 = _T_2327 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_285 = _T_2328 | vArrayWire_31_2; // @[Reg.scala 28:19]
  wire  _T_2340 = selArrayWire_31 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2341 = _T_2294 & _T_2340; // @[Cache.scala 114:85]
  wire  _T_2342 = _T_2341 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_287 = _T_2342 | vArrayWire_31_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2353 = selArrayWire_32 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2355 = io_cacheOut_r_last_i & _T_191; // @[Cache.scala 111:28]
  wire  _T_2359 = selArrayWire_32 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2360 = _T_2355 & _T_2359; // @[Cache.scala 114:85]
  wire  _T_2361 = _T_2360 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_290 = _T_2361 | vArrayWire_32_0; // @[Reg.scala 28:19]
  wire  _T_2373 = selArrayWire_32 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2374 = _T_2355 & _T_2373; // @[Cache.scala 114:85]
  wire  _T_2375 = _T_2374 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_292 = _T_2375 | vArrayWire_32_1; // @[Reg.scala 28:19]
  wire  _T_2387 = selArrayWire_32 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2388 = _T_2355 & _T_2387; // @[Cache.scala 114:85]
  wire  _T_2389 = _T_2388 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_294 = _T_2389 | vArrayWire_32_2; // @[Reg.scala 28:19]
  wire  _T_2401 = selArrayWire_32 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2402 = _T_2355 & _T_2401; // @[Cache.scala 114:85]
  wire  _T_2403 = _T_2402 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_296 = _T_2403 | vArrayWire_32_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2414 = selArrayWire_33 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2416 = io_cacheOut_r_last_i & _T_193; // @[Cache.scala 111:28]
  wire  _T_2420 = selArrayWire_33 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2421 = _T_2416 & _T_2420; // @[Cache.scala 114:85]
  wire  _T_2422 = _T_2421 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_299 = _T_2422 | vArrayWire_33_0; // @[Reg.scala 28:19]
  wire  _T_2434 = selArrayWire_33 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2435 = _T_2416 & _T_2434; // @[Cache.scala 114:85]
  wire  _T_2436 = _T_2435 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_301 = _T_2436 | vArrayWire_33_1; // @[Reg.scala 28:19]
  wire  _T_2448 = selArrayWire_33 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2449 = _T_2416 & _T_2448; // @[Cache.scala 114:85]
  wire  _T_2450 = _T_2449 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_303 = _T_2450 | vArrayWire_33_2; // @[Reg.scala 28:19]
  wire  _T_2462 = selArrayWire_33 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2463 = _T_2416 & _T_2462; // @[Cache.scala 114:85]
  wire  _T_2464 = _T_2463 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_305 = _T_2464 | vArrayWire_33_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2475 = selArrayWire_34 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2477 = io_cacheOut_r_last_i & _T_195; // @[Cache.scala 111:28]
  wire  _T_2481 = selArrayWire_34 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2482 = _T_2477 & _T_2481; // @[Cache.scala 114:85]
  wire  _T_2483 = _T_2482 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_308 = _T_2483 | vArrayWire_34_0; // @[Reg.scala 28:19]
  wire  _T_2495 = selArrayWire_34 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2496 = _T_2477 & _T_2495; // @[Cache.scala 114:85]
  wire  _T_2497 = _T_2496 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_310 = _T_2497 | vArrayWire_34_1; // @[Reg.scala 28:19]
  wire  _T_2509 = selArrayWire_34 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2510 = _T_2477 & _T_2509; // @[Cache.scala 114:85]
  wire  _T_2511 = _T_2510 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_312 = _T_2511 | vArrayWire_34_2; // @[Reg.scala 28:19]
  wire  _T_2523 = selArrayWire_34 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2524 = _T_2477 & _T_2523; // @[Cache.scala 114:85]
  wire  _T_2525 = _T_2524 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_314 = _T_2525 | vArrayWire_34_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2536 = selArrayWire_35 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2538 = io_cacheOut_r_last_i & _T_197; // @[Cache.scala 111:28]
  wire  _T_2542 = selArrayWire_35 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2543 = _T_2538 & _T_2542; // @[Cache.scala 114:85]
  wire  _T_2544 = _T_2543 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_317 = _T_2544 | vArrayWire_35_0; // @[Reg.scala 28:19]
  wire  _T_2556 = selArrayWire_35 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2557 = _T_2538 & _T_2556; // @[Cache.scala 114:85]
  wire  _T_2558 = _T_2557 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_319 = _T_2558 | vArrayWire_35_1; // @[Reg.scala 28:19]
  wire  _T_2570 = selArrayWire_35 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2571 = _T_2538 & _T_2570; // @[Cache.scala 114:85]
  wire  _T_2572 = _T_2571 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_321 = _T_2572 | vArrayWire_35_2; // @[Reg.scala 28:19]
  wire  _T_2584 = selArrayWire_35 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2585 = _T_2538 & _T_2584; // @[Cache.scala 114:85]
  wire  _T_2586 = _T_2585 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_323 = _T_2586 | vArrayWire_35_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2597 = selArrayWire_36 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2599 = io_cacheOut_r_last_i & _T_199; // @[Cache.scala 111:28]
  wire  _T_2603 = selArrayWire_36 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2604 = _T_2599 & _T_2603; // @[Cache.scala 114:85]
  wire  _T_2605 = _T_2604 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_326 = _T_2605 | vArrayWire_36_0; // @[Reg.scala 28:19]
  wire  _T_2617 = selArrayWire_36 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2618 = _T_2599 & _T_2617; // @[Cache.scala 114:85]
  wire  _T_2619 = _T_2618 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_328 = _T_2619 | vArrayWire_36_1; // @[Reg.scala 28:19]
  wire  _T_2631 = selArrayWire_36 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2632 = _T_2599 & _T_2631; // @[Cache.scala 114:85]
  wire  _T_2633 = _T_2632 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_330 = _T_2633 | vArrayWire_36_2; // @[Reg.scala 28:19]
  wire  _T_2645 = selArrayWire_36 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2646 = _T_2599 & _T_2645; // @[Cache.scala 114:85]
  wire  _T_2647 = _T_2646 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_332 = _T_2647 | vArrayWire_36_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2658 = selArrayWire_37 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2660 = io_cacheOut_r_last_i & _T_201; // @[Cache.scala 111:28]
  wire  _T_2664 = selArrayWire_37 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2665 = _T_2660 & _T_2664; // @[Cache.scala 114:85]
  wire  _T_2666 = _T_2665 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_335 = _T_2666 | vArrayWire_37_0; // @[Reg.scala 28:19]
  wire  _T_2678 = selArrayWire_37 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2679 = _T_2660 & _T_2678; // @[Cache.scala 114:85]
  wire  _T_2680 = _T_2679 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_337 = _T_2680 | vArrayWire_37_1; // @[Reg.scala 28:19]
  wire  _T_2692 = selArrayWire_37 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2693 = _T_2660 & _T_2692; // @[Cache.scala 114:85]
  wire  _T_2694 = _T_2693 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_339 = _T_2694 | vArrayWire_37_2; // @[Reg.scala 28:19]
  wire  _T_2706 = selArrayWire_37 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2707 = _T_2660 & _T_2706; // @[Cache.scala 114:85]
  wire  _T_2708 = _T_2707 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_341 = _T_2708 | vArrayWire_37_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2719 = selArrayWire_38 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2721 = io_cacheOut_r_last_i & _T_203; // @[Cache.scala 111:28]
  wire  _T_2725 = selArrayWire_38 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2726 = _T_2721 & _T_2725; // @[Cache.scala 114:85]
  wire  _T_2727 = _T_2726 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_344 = _T_2727 | vArrayWire_38_0; // @[Reg.scala 28:19]
  wire  _T_2739 = selArrayWire_38 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2740 = _T_2721 & _T_2739; // @[Cache.scala 114:85]
  wire  _T_2741 = _T_2740 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_346 = _T_2741 | vArrayWire_38_1; // @[Reg.scala 28:19]
  wire  _T_2753 = selArrayWire_38 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2754 = _T_2721 & _T_2753; // @[Cache.scala 114:85]
  wire  _T_2755 = _T_2754 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_348 = _T_2755 | vArrayWire_38_2; // @[Reg.scala 28:19]
  wire  _T_2767 = selArrayWire_38 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2768 = _T_2721 & _T_2767; // @[Cache.scala 114:85]
  wire  _T_2769 = _T_2768 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_350 = _T_2769 | vArrayWire_38_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2780 = selArrayWire_39 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2782 = io_cacheOut_r_last_i & _T_205; // @[Cache.scala 111:28]
  wire  _T_2786 = selArrayWire_39 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2787 = _T_2782 & _T_2786; // @[Cache.scala 114:85]
  wire  _T_2788 = _T_2787 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_353 = _T_2788 | vArrayWire_39_0; // @[Reg.scala 28:19]
  wire  _T_2800 = selArrayWire_39 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2801 = _T_2782 & _T_2800; // @[Cache.scala 114:85]
  wire  _T_2802 = _T_2801 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_355 = _T_2802 | vArrayWire_39_1; // @[Reg.scala 28:19]
  wire  _T_2814 = selArrayWire_39 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2815 = _T_2782 & _T_2814; // @[Cache.scala 114:85]
  wire  _T_2816 = _T_2815 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_357 = _T_2816 | vArrayWire_39_2; // @[Reg.scala 28:19]
  wire  _T_2828 = selArrayWire_39 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2829 = _T_2782 & _T_2828; // @[Cache.scala 114:85]
  wire  _T_2830 = _T_2829 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_359 = _T_2830 | vArrayWire_39_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2841 = selArrayWire_40 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2843 = io_cacheOut_r_last_i & _T_207; // @[Cache.scala 111:28]
  wire  _T_2847 = selArrayWire_40 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2848 = _T_2843 & _T_2847; // @[Cache.scala 114:85]
  wire  _T_2849 = _T_2848 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_362 = _T_2849 | vArrayWire_40_0; // @[Reg.scala 28:19]
  wire  _T_2861 = selArrayWire_40 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2862 = _T_2843 & _T_2861; // @[Cache.scala 114:85]
  wire  _T_2863 = _T_2862 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_364 = _T_2863 | vArrayWire_40_1; // @[Reg.scala 28:19]
  wire  _T_2875 = selArrayWire_40 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2876 = _T_2843 & _T_2875; // @[Cache.scala 114:85]
  wire  _T_2877 = _T_2876 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_366 = _T_2877 | vArrayWire_40_2; // @[Reg.scala 28:19]
  wire  _T_2889 = selArrayWire_40 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2890 = _T_2843 & _T_2889; // @[Cache.scala 114:85]
  wire  _T_2891 = _T_2890 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_368 = _T_2891 | vArrayWire_40_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2902 = selArrayWire_41 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2904 = io_cacheOut_r_last_i & _T_209; // @[Cache.scala 111:28]
  wire  _T_2908 = selArrayWire_41 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2909 = _T_2904 & _T_2908; // @[Cache.scala 114:85]
  wire  _T_2910 = _T_2909 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_371 = _T_2910 | vArrayWire_41_0; // @[Reg.scala 28:19]
  wire  _T_2922 = selArrayWire_41 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2923 = _T_2904 & _T_2922; // @[Cache.scala 114:85]
  wire  _T_2924 = _T_2923 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_373 = _T_2924 | vArrayWire_41_1; // @[Reg.scala 28:19]
  wire  _T_2936 = selArrayWire_41 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2937 = _T_2904 & _T_2936; // @[Cache.scala 114:85]
  wire  _T_2938 = _T_2937 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_375 = _T_2938 | vArrayWire_41_2; // @[Reg.scala 28:19]
  wire  _T_2950 = selArrayWire_41 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_2951 = _T_2904 & _T_2950; // @[Cache.scala 114:85]
  wire  _T_2952 = _T_2951 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_377 = _T_2952 | vArrayWire_41_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2963 = selArrayWire_42 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_2965 = io_cacheOut_r_last_i & _T_211; // @[Cache.scala 111:28]
  wire  _T_2969 = selArrayWire_42 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_2970 = _T_2965 & _T_2969; // @[Cache.scala 114:85]
  wire  _T_2971 = _T_2970 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_380 = _T_2971 | vArrayWire_42_0; // @[Reg.scala 28:19]
  wire  _T_2983 = selArrayWire_42 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_2984 = _T_2965 & _T_2983; // @[Cache.scala 114:85]
  wire  _T_2985 = _T_2984 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_382 = _T_2985 | vArrayWire_42_1; // @[Reg.scala 28:19]
  wire  _T_2997 = selArrayWire_42 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_2998 = _T_2965 & _T_2997; // @[Cache.scala 114:85]
  wire  _T_2999 = _T_2998 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_384 = _T_2999 | vArrayWire_42_2; // @[Reg.scala 28:19]
  wire  _T_3011 = selArrayWire_42 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3012 = _T_2965 & _T_3011; // @[Cache.scala 114:85]
  wire  _T_3013 = _T_3012 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_386 = _T_3013 | vArrayWire_42_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3024 = selArrayWire_43 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3026 = io_cacheOut_r_last_i & _T_213; // @[Cache.scala 111:28]
  wire  _T_3030 = selArrayWire_43 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3031 = _T_3026 & _T_3030; // @[Cache.scala 114:85]
  wire  _T_3032 = _T_3031 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_389 = _T_3032 | vArrayWire_43_0; // @[Reg.scala 28:19]
  wire  _T_3044 = selArrayWire_43 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3045 = _T_3026 & _T_3044; // @[Cache.scala 114:85]
  wire  _T_3046 = _T_3045 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_391 = _T_3046 | vArrayWire_43_1; // @[Reg.scala 28:19]
  wire  _T_3058 = selArrayWire_43 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3059 = _T_3026 & _T_3058; // @[Cache.scala 114:85]
  wire  _T_3060 = _T_3059 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_393 = _T_3060 | vArrayWire_43_2; // @[Reg.scala 28:19]
  wire  _T_3072 = selArrayWire_43 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3073 = _T_3026 & _T_3072; // @[Cache.scala 114:85]
  wire  _T_3074 = _T_3073 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_395 = _T_3074 | vArrayWire_43_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3085 = selArrayWire_44 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3087 = io_cacheOut_r_last_i & _T_215; // @[Cache.scala 111:28]
  wire  _T_3091 = selArrayWire_44 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3092 = _T_3087 & _T_3091; // @[Cache.scala 114:85]
  wire  _T_3093 = _T_3092 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_398 = _T_3093 | vArrayWire_44_0; // @[Reg.scala 28:19]
  wire  _T_3105 = selArrayWire_44 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3106 = _T_3087 & _T_3105; // @[Cache.scala 114:85]
  wire  _T_3107 = _T_3106 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_400 = _T_3107 | vArrayWire_44_1; // @[Reg.scala 28:19]
  wire  _T_3119 = selArrayWire_44 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3120 = _T_3087 & _T_3119; // @[Cache.scala 114:85]
  wire  _T_3121 = _T_3120 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_402 = _T_3121 | vArrayWire_44_2; // @[Reg.scala 28:19]
  wire  _T_3133 = selArrayWire_44 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3134 = _T_3087 & _T_3133; // @[Cache.scala 114:85]
  wire  _T_3135 = _T_3134 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_404 = _T_3135 | vArrayWire_44_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3146 = selArrayWire_45 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3148 = io_cacheOut_r_last_i & _T_217; // @[Cache.scala 111:28]
  wire  _T_3152 = selArrayWire_45 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3153 = _T_3148 & _T_3152; // @[Cache.scala 114:85]
  wire  _T_3154 = _T_3153 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_407 = _T_3154 | vArrayWire_45_0; // @[Reg.scala 28:19]
  wire  _T_3166 = selArrayWire_45 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3167 = _T_3148 & _T_3166; // @[Cache.scala 114:85]
  wire  _T_3168 = _T_3167 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_409 = _T_3168 | vArrayWire_45_1; // @[Reg.scala 28:19]
  wire  _T_3180 = selArrayWire_45 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3181 = _T_3148 & _T_3180; // @[Cache.scala 114:85]
  wire  _T_3182 = _T_3181 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_411 = _T_3182 | vArrayWire_45_2; // @[Reg.scala 28:19]
  wire  _T_3194 = selArrayWire_45 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3195 = _T_3148 & _T_3194; // @[Cache.scala 114:85]
  wire  _T_3196 = _T_3195 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_413 = _T_3196 | vArrayWire_45_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3207 = selArrayWire_46 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3209 = io_cacheOut_r_last_i & _T_219; // @[Cache.scala 111:28]
  wire  _T_3213 = selArrayWire_46 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3214 = _T_3209 & _T_3213; // @[Cache.scala 114:85]
  wire  _T_3215 = _T_3214 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_416 = _T_3215 | vArrayWire_46_0; // @[Reg.scala 28:19]
  wire  _T_3227 = selArrayWire_46 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3228 = _T_3209 & _T_3227; // @[Cache.scala 114:85]
  wire  _T_3229 = _T_3228 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_418 = _T_3229 | vArrayWire_46_1; // @[Reg.scala 28:19]
  wire  _T_3241 = selArrayWire_46 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3242 = _T_3209 & _T_3241; // @[Cache.scala 114:85]
  wire  _T_3243 = _T_3242 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_420 = _T_3243 | vArrayWire_46_2; // @[Reg.scala 28:19]
  wire  _T_3255 = selArrayWire_46 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3256 = _T_3209 & _T_3255; // @[Cache.scala 114:85]
  wire  _T_3257 = _T_3256 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_422 = _T_3257 | vArrayWire_46_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3268 = selArrayWire_47 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3270 = io_cacheOut_r_last_i & _T_221; // @[Cache.scala 111:28]
  wire  _T_3274 = selArrayWire_47 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3275 = _T_3270 & _T_3274; // @[Cache.scala 114:85]
  wire  _T_3276 = _T_3275 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_425 = _T_3276 | vArrayWire_47_0; // @[Reg.scala 28:19]
  wire  _T_3288 = selArrayWire_47 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3289 = _T_3270 & _T_3288; // @[Cache.scala 114:85]
  wire  _T_3290 = _T_3289 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_427 = _T_3290 | vArrayWire_47_1; // @[Reg.scala 28:19]
  wire  _T_3302 = selArrayWire_47 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3303 = _T_3270 & _T_3302; // @[Cache.scala 114:85]
  wire  _T_3304 = _T_3303 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_429 = _T_3304 | vArrayWire_47_2; // @[Reg.scala 28:19]
  wire  _T_3316 = selArrayWire_47 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3317 = _T_3270 & _T_3316; // @[Cache.scala 114:85]
  wire  _T_3318 = _T_3317 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_431 = _T_3318 | vArrayWire_47_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3329 = selArrayWire_48 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3331 = io_cacheOut_r_last_i & _T_223; // @[Cache.scala 111:28]
  wire  _T_3335 = selArrayWire_48 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3336 = _T_3331 & _T_3335; // @[Cache.scala 114:85]
  wire  _T_3337 = _T_3336 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_434 = _T_3337 | vArrayWire_48_0; // @[Reg.scala 28:19]
  wire  _T_3349 = selArrayWire_48 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3350 = _T_3331 & _T_3349; // @[Cache.scala 114:85]
  wire  _T_3351 = _T_3350 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_436 = _T_3351 | vArrayWire_48_1; // @[Reg.scala 28:19]
  wire  _T_3363 = selArrayWire_48 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3364 = _T_3331 & _T_3363; // @[Cache.scala 114:85]
  wire  _T_3365 = _T_3364 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_438 = _T_3365 | vArrayWire_48_2; // @[Reg.scala 28:19]
  wire  _T_3377 = selArrayWire_48 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3378 = _T_3331 & _T_3377; // @[Cache.scala 114:85]
  wire  _T_3379 = _T_3378 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_440 = _T_3379 | vArrayWire_48_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3390 = selArrayWire_49 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3392 = io_cacheOut_r_last_i & _T_225; // @[Cache.scala 111:28]
  wire  _T_3396 = selArrayWire_49 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3397 = _T_3392 & _T_3396; // @[Cache.scala 114:85]
  wire  _T_3398 = _T_3397 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_443 = _T_3398 | vArrayWire_49_0; // @[Reg.scala 28:19]
  wire  _T_3410 = selArrayWire_49 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3411 = _T_3392 & _T_3410; // @[Cache.scala 114:85]
  wire  _T_3412 = _T_3411 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_445 = _T_3412 | vArrayWire_49_1; // @[Reg.scala 28:19]
  wire  _T_3424 = selArrayWire_49 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3425 = _T_3392 & _T_3424; // @[Cache.scala 114:85]
  wire  _T_3426 = _T_3425 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_447 = _T_3426 | vArrayWire_49_2; // @[Reg.scala 28:19]
  wire  _T_3438 = selArrayWire_49 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3439 = _T_3392 & _T_3438; // @[Cache.scala 114:85]
  wire  _T_3440 = _T_3439 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_449 = _T_3440 | vArrayWire_49_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3451 = selArrayWire_50 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3453 = io_cacheOut_r_last_i & _T_227; // @[Cache.scala 111:28]
  wire  _T_3457 = selArrayWire_50 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3458 = _T_3453 & _T_3457; // @[Cache.scala 114:85]
  wire  _T_3459 = _T_3458 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_452 = _T_3459 | vArrayWire_50_0; // @[Reg.scala 28:19]
  wire  _T_3471 = selArrayWire_50 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3472 = _T_3453 & _T_3471; // @[Cache.scala 114:85]
  wire  _T_3473 = _T_3472 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_454 = _T_3473 | vArrayWire_50_1; // @[Reg.scala 28:19]
  wire  _T_3485 = selArrayWire_50 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3486 = _T_3453 & _T_3485; // @[Cache.scala 114:85]
  wire  _T_3487 = _T_3486 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_456 = _T_3487 | vArrayWire_50_2; // @[Reg.scala 28:19]
  wire  _T_3499 = selArrayWire_50 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3500 = _T_3453 & _T_3499; // @[Cache.scala 114:85]
  wire  _T_3501 = _T_3500 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_458 = _T_3501 | vArrayWire_50_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3512 = selArrayWire_51 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3514 = io_cacheOut_r_last_i & _T_229; // @[Cache.scala 111:28]
  wire  _T_3518 = selArrayWire_51 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3519 = _T_3514 & _T_3518; // @[Cache.scala 114:85]
  wire  _T_3520 = _T_3519 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_461 = _T_3520 | vArrayWire_51_0; // @[Reg.scala 28:19]
  wire  _T_3532 = selArrayWire_51 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3533 = _T_3514 & _T_3532; // @[Cache.scala 114:85]
  wire  _T_3534 = _T_3533 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_463 = _T_3534 | vArrayWire_51_1; // @[Reg.scala 28:19]
  wire  _T_3546 = selArrayWire_51 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3547 = _T_3514 & _T_3546; // @[Cache.scala 114:85]
  wire  _T_3548 = _T_3547 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_465 = _T_3548 | vArrayWire_51_2; // @[Reg.scala 28:19]
  wire  _T_3560 = selArrayWire_51 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3561 = _T_3514 & _T_3560; // @[Cache.scala 114:85]
  wire  _T_3562 = _T_3561 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_467 = _T_3562 | vArrayWire_51_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3573 = selArrayWire_52 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3575 = io_cacheOut_r_last_i & _T_231; // @[Cache.scala 111:28]
  wire  _T_3579 = selArrayWire_52 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3580 = _T_3575 & _T_3579; // @[Cache.scala 114:85]
  wire  _T_3581 = _T_3580 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_470 = _T_3581 | vArrayWire_52_0; // @[Reg.scala 28:19]
  wire  _T_3593 = selArrayWire_52 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3594 = _T_3575 & _T_3593; // @[Cache.scala 114:85]
  wire  _T_3595 = _T_3594 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_472 = _T_3595 | vArrayWire_52_1; // @[Reg.scala 28:19]
  wire  _T_3607 = selArrayWire_52 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3608 = _T_3575 & _T_3607; // @[Cache.scala 114:85]
  wire  _T_3609 = _T_3608 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_474 = _T_3609 | vArrayWire_52_2; // @[Reg.scala 28:19]
  wire  _T_3621 = selArrayWire_52 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3622 = _T_3575 & _T_3621; // @[Cache.scala 114:85]
  wire  _T_3623 = _T_3622 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_476 = _T_3623 | vArrayWire_52_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3634 = selArrayWire_53 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3636 = io_cacheOut_r_last_i & _T_233; // @[Cache.scala 111:28]
  wire  _T_3640 = selArrayWire_53 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3641 = _T_3636 & _T_3640; // @[Cache.scala 114:85]
  wire  _T_3642 = _T_3641 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_479 = _T_3642 | vArrayWire_53_0; // @[Reg.scala 28:19]
  wire  _T_3654 = selArrayWire_53 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3655 = _T_3636 & _T_3654; // @[Cache.scala 114:85]
  wire  _T_3656 = _T_3655 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_481 = _T_3656 | vArrayWire_53_1; // @[Reg.scala 28:19]
  wire  _T_3668 = selArrayWire_53 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3669 = _T_3636 & _T_3668; // @[Cache.scala 114:85]
  wire  _T_3670 = _T_3669 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_483 = _T_3670 | vArrayWire_53_2; // @[Reg.scala 28:19]
  wire  _T_3682 = selArrayWire_53 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3683 = _T_3636 & _T_3682; // @[Cache.scala 114:85]
  wire  _T_3684 = _T_3683 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_485 = _T_3684 | vArrayWire_53_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3695 = selArrayWire_54 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3697 = io_cacheOut_r_last_i & _T_235; // @[Cache.scala 111:28]
  wire  _T_3701 = selArrayWire_54 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3702 = _T_3697 & _T_3701; // @[Cache.scala 114:85]
  wire  _T_3703 = _T_3702 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_488 = _T_3703 | vArrayWire_54_0; // @[Reg.scala 28:19]
  wire  _T_3715 = selArrayWire_54 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3716 = _T_3697 & _T_3715; // @[Cache.scala 114:85]
  wire  _T_3717 = _T_3716 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_490 = _T_3717 | vArrayWire_54_1; // @[Reg.scala 28:19]
  wire  _T_3729 = selArrayWire_54 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3730 = _T_3697 & _T_3729; // @[Cache.scala 114:85]
  wire  _T_3731 = _T_3730 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_492 = _T_3731 | vArrayWire_54_2; // @[Reg.scala 28:19]
  wire  _T_3743 = selArrayWire_54 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3744 = _T_3697 & _T_3743; // @[Cache.scala 114:85]
  wire  _T_3745 = _T_3744 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_494 = _T_3745 | vArrayWire_54_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3756 = selArrayWire_55 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3758 = io_cacheOut_r_last_i & _T_237; // @[Cache.scala 111:28]
  wire  _T_3762 = selArrayWire_55 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3763 = _T_3758 & _T_3762; // @[Cache.scala 114:85]
  wire  _T_3764 = _T_3763 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_497 = _T_3764 | vArrayWire_55_0; // @[Reg.scala 28:19]
  wire  _T_3776 = selArrayWire_55 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3777 = _T_3758 & _T_3776; // @[Cache.scala 114:85]
  wire  _T_3778 = _T_3777 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_499 = _T_3778 | vArrayWire_55_1; // @[Reg.scala 28:19]
  wire  _T_3790 = selArrayWire_55 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3791 = _T_3758 & _T_3790; // @[Cache.scala 114:85]
  wire  _T_3792 = _T_3791 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_501 = _T_3792 | vArrayWire_55_2; // @[Reg.scala 28:19]
  wire  _T_3804 = selArrayWire_55 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3805 = _T_3758 & _T_3804; // @[Cache.scala 114:85]
  wire  _T_3806 = _T_3805 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_503 = _T_3806 | vArrayWire_55_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3817 = selArrayWire_56 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3819 = io_cacheOut_r_last_i & _T_239; // @[Cache.scala 111:28]
  wire  _T_3823 = selArrayWire_56 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3824 = _T_3819 & _T_3823; // @[Cache.scala 114:85]
  wire  _T_3825 = _T_3824 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_506 = _T_3825 | vArrayWire_56_0; // @[Reg.scala 28:19]
  wire  _T_3837 = selArrayWire_56 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3838 = _T_3819 & _T_3837; // @[Cache.scala 114:85]
  wire  _T_3839 = _T_3838 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_508 = _T_3839 | vArrayWire_56_1; // @[Reg.scala 28:19]
  wire  _T_3851 = selArrayWire_56 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3852 = _T_3819 & _T_3851; // @[Cache.scala 114:85]
  wire  _T_3853 = _T_3852 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_510 = _T_3853 | vArrayWire_56_2; // @[Reg.scala 28:19]
  wire  _T_3865 = selArrayWire_56 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3866 = _T_3819 & _T_3865; // @[Cache.scala 114:85]
  wire  _T_3867 = _T_3866 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_512 = _T_3867 | vArrayWire_56_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3878 = selArrayWire_57 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3880 = io_cacheOut_r_last_i & _T_241; // @[Cache.scala 111:28]
  wire  _T_3884 = selArrayWire_57 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3885 = _T_3880 & _T_3884; // @[Cache.scala 114:85]
  wire  _T_3886 = _T_3885 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_515 = _T_3886 | vArrayWire_57_0; // @[Reg.scala 28:19]
  wire  _T_3898 = selArrayWire_57 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3899 = _T_3880 & _T_3898; // @[Cache.scala 114:85]
  wire  _T_3900 = _T_3899 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_517 = _T_3900 | vArrayWire_57_1; // @[Reg.scala 28:19]
  wire  _T_3912 = selArrayWire_57 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3913 = _T_3880 & _T_3912; // @[Cache.scala 114:85]
  wire  _T_3914 = _T_3913 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_519 = _T_3914 | vArrayWire_57_2; // @[Reg.scala 28:19]
  wire  _T_3926 = selArrayWire_57 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3927 = _T_3880 & _T_3926; // @[Cache.scala 114:85]
  wire  _T_3928 = _T_3927 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_521 = _T_3928 | vArrayWire_57_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3939 = selArrayWire_58 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_3941 = io_cacheOut_r_last_i & _T_243; // @[Cache.scala 111:28]
  wire  _T_3945 = selArrayWire_58 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_3946 = _T_3941 & _T_3945; // @[Cache.scala 114:85]
  wire  _T_3947 = _T_3946 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_524 = _T_3947 | vArrayWire_58_0; // @[Reg.scala 28:19]
  wire  _T_3959 = selArrayWire_58 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_3960 = _T_3941 & _T_3959; // @[Cache.scala 114:85]
  wire  _T_3961 = _T_3960 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_526 = _T_3961 | vArrayWire_58_1; // @[Reg.scala 28:19]
  wire  _T_3973 = selArrayWire_58 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_3974 = _T_3941 & _T_3973; // @[Cache.scala 114:85]
  wire  _T_3975 = _T_3974 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_528 = _T_3975 | vArrayWire_58_2; // @[Reg.scala 28:19]
  wire  _T_3987 = selArrayWire_58 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_3988 = _T_3941 & _T_3987; // @[Cache.scala 114:85]
  wire  _T_3989 = _T_3988 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_530 = _T_3989 | vArrayWire_58_3; // @[Reg.scala 28:19]
  wire [1:0] _T_4000 = selArrayWire_59 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_4002 = io_cacheOut_r_last_i & _T_245; // @[Cache.scala 111:28]
  wire  _T_4006 = selArrayWire_59 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_4007 = _T_4002 & _T_4006; // @[Cache.scala 114:85]
  wire  _T_4008 = _T_4007 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_533 = _T_4008 | vArrayWire_59_0; // @[Reg.scala 28:19]
  wire  _T_4020 = selArrayWire_59 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_4021 = _T_4002 & _T_4020; // @[Cache.scala 114:85]
  wire  _T_4022 = _T_4021 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_535 = _T_4022 | vArrayWire_59_1; // @[Reg.scala 28:19]
  wire  _T_4034 = selArrayWire_59 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_4035 = _T_4002 & _T_4034; // @[Cache.scala 114:85]
  wire  _T_4036 = _T_4035 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_537 = _T_4036 | vArrayWire_59_2; // @[Reg.scala 28:19]
  wire  _T_4048 = selArrayWire_59 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_4049 = _T_4002 & _T_4048; // @[Cache.scala 114:85]
  wire  _T_4050 = _T_4049 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_539 = _T_4050 | vArrayWire_59_3; // @[Reg.scala 28:19]
  wire [1:0] _T_4061 = selArrayWire_60 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_4063 = io_cacheOut_r_last_i & _T_247; // @[Cache.scala 111:28]
  wire  _T_4067 = selArrayWire_60 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_4068 = _T_4063 & _T_4067; // @[Cache.scala 114:85]
  wire  _T_4069 = _T_4068 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_542 = _T_4069 | vArrayWire_60_0; // @[Reg.scala 28:19]
  wire  _T_4081 = selArrayWire_60 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_4082 = _T_4063 & _T_4081; // @[Cache.scala 114:85]
  wire  _T_4083 = _T_4082 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_544 = _T_4083 | vArrayWire_60_1; // @[Reg.scala 28:19]
  wire  _T_4095 = selArrayWire_60 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_4096 = _T_4063 & _T_4095; // @[Cache.scala 114:85]
  wire  _T_4097 = _T_4096 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_546 = _T_4097 | vArrayWire_60_2; // @[Reg.scala 28:19]
  wire  _T_4109 = selArrayWire_60 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_4110 = _T_4063 & _T_4109; // @[Cache.scala 114:85]
  wire  _T_4111 = _T_4110 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_548 = _T_4111 | vArrayWire_60_3; // @[Reg.scala 28:19]
  wire [1:0] _T_4122 = selArrayWire_61 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_4124 = io_cacheOut_r_last_i & _T_249; // @[Cache.scala 111:28]
  wire  _T_4128 = selArrayWire_61 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_4129 = _T_4124 & _T_4128; // @[Cache.scala 114:85]
  wire  _T_4130 = _T_4129 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_551 = _T_4130 | vArrayWire_61_0; // @[Reg.scala 28:19]
  wire  _T_4142 = selArrayWire_61 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_4143 = _T_4124 & _T_4142; // @[Cache.scala 114:85]
  wire  _T_4144 = _T_4143 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_553 = _T_4144 | vArrayWire_61_1; // @[Reg.scala 28:19]
  wire  _T_4156 = selArrayWire_61 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_4157 = _T_4124 & _T_4156; // @[Cache.scala 114:85]
  wire  _T_4158 = _T_4157 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_555 = _T_4158 | vArrayWire_61_2; // @[Reg.scala 28:19]
  wire  _T_4170 = selArrayWire_61 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_4171 = _T_4124 & _T_4170; // @[Cache.scala 114:85]
  wire  _T_4172 = _T_4171 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_557 = _T_4172 | vArrayWire_61_3; // @[Reg.scala 28:19]
  wire [1:0] _T_4183 = selArrayWire_62 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_4185 = io_cacheOut_r_last_i & _T_251; // @[Cache.scala 111:28]
  wire  _T_4189 = selArrayWire_62 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_4190 = _T_4185 & _T_4189; // @[Cache.scala 114:85]
  wire  _T_4191 = _T_4190 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_560 = _T_4191 | vArrayWire_62_0; // @[Reg.scala 28:19]
  wire  _T_4203 = selArrayWire_62 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_4204 = _T_4185 & _T_4203; // @[Cache.scala 114:85]
  wire  _T_4205 = _T_4204 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_562 = _T_4205 | vArrayWire_62_1; // @[Reg.scala 28:19]
  wire  _T_4217 = selArrayWire_62 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_4218 = _T_4185 & _T_4217; // @[Cache.scala 114:85]
  wire  _T_4219 = _T_4218 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_564 = _T_4219 | vArrayWire_62_2; // @[Reg.scala 28:19]
  wire  _T_4231 = selArrayWire_62 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_4232 = _T_4185 & _T_4231; // @[Cache.scala 114:85]
  wire  _T_4233 = _T_4232 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_566 = _T_4233 | vArrayWire_62_3; // @[Reg.scala 28:19]
  wire [1:0] _T_4244 = selArrayWire_63 + 2'h1; // @[Cache.scala 109:23]
  wire  _T_4246 = io_cacheOut_r_last_i & _T_253; // @[Cache.scala 111:28]
  wire  _T_4250 = selArrayWire_63 == 2'h0; // @[Cache.scala 114:104]
  wire  _T_4251 = _T_4246 & _T_4250; // @[Cache.scala 114:85]
  wire  _T_4252 = _T_4251 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_569 = _T_4252 | vArrayWire_63_0; // @[Reg.scala 28:19]
  wire  _T_4264 = selArrayWire_63 == 2'h1; // @[Cache.scala 114:104]
  wire  _T_4265 = _T_4246 & _T_4264; // @[Cache.scala 114:85]
  wire  _T_4266 = _T_4265 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_571 = _T_4266 | vArrayWire_63_1; // @[Reg.scala 28:19]
  wire  _T_4278 = selArrayWire_63 == 2'h2; // @[Cache.scala 114:104]
  wire  _T_4279 = _T_4246 & _T_4278; // @[Cache.scala 114:85]
  wire  _T_4280 = _T_4279 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_573 = _T_4280 | vArrayWire_63_2; // @[Reg.scala 28:19]
  wire  _T_4292 = selArrayWire_63 == 2'h3; // @[Cache.scala 114:104]
  wire  _T_4293 = _T_4246 & _T_4292; // @[Cache.scala 114:85]
  wire  _T_4294 = _T_4293 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_575 = _T_4294 | vArrayWire_63_3; // @[Reg.scala 28:19]
  wire  _T_4357 = cacheState & io_cacheOut_r_valid_i; // @[Cache.scala 147:26]
  wire  _T_4358 = 2'h0 == sramSel; // @[Cache.scala 147:61]
  wire  _T_4359 = _T_4357 & _T_4358; // @[Cache.scala 147:52]
  wire [127:0] _T_4365 = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_4366 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 29:58]
  wire  _T_4376 = 2'h1 == sramSel; // @[Cache.scala 147:61]
  wire  _T_4377 = _T_4357 & _T_4376; // @[Cache.scala 147:52]
  wire  _T_4394 = 2'h2 == sramSel; // @[Cache.scala 147:61]
  wire  _T_4395 = _T_4357 & _T_4394; // @[Cache.scala 147:52]
  wire  _T_4412 = 2'h3 == sramSel; // @[Cache.scala 147:61]
  wire  _T_4413 = _T_4357 & _T_4412; // @[Cache.scala 147:52]
  assign io_cacheOut_ar_valid_o = cacheState; // @[Cache.scala 105:26]
  assign io_cacheOut_ar_addr_o = {io_cacheIn_addr[31:4],4'h0}; // @[Cache.scala 104:25]
  assign io_cacheOut_ar_len_o = {{7'd0}, cacheState}; // @[Cache.scala 103:24]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 139:24]
  assign io_cacheIn_ready = isIdle & hit; // @[Cache.scala 155:20]
  assign io_cacheIn_data_read = offset[3] ? waysel[127:64] : waysel[63:0]; // @[Cache.scala 92:24]
  assign io_SRAMIO_0_cen = ~_T_4359; // @[Cache.scala 147:13]
  assign io_SRAMIO_0_wen = ~_T_4359; // @[Cache.scala 149:13]
  assign io_SRAMIO_0_wdata = io_cacheOut_r_last_i ? _T_4365 : _T_4366; // @[Cache.scala 150:15]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 148:14]
  assign io_SRAMIO_0_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:15]
  assign io_SRAMIO_1_cen = ~_T_4377; // @[Cache.scala 147:13]
  assign io_SRAMIO_1_wen = ~_T_4377; // @[Cache.scala 149:13]
  assign io_SRAMIO_1_wdata = io_cacheOut_r_last_i ? _T_4365 : _T_4366; // @[Cache.scala 150:15]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 148:14]
  assign io_SRAMIO_1_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:15]
  assign io_SRAMIO_2_cen = ~_T_4395; // @[Cache.scala 147:13]
  assign io_SRAMIO_2_wen = ~_T_4395; // @[Cache.scala 149:13]
  assign io_SRAMIO_2_wdata = io_cacheOut_r_last_i ? _T_4365 : _T_4366; // @[Cache.scala 150:15]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 148:14]
  assign io_SRAMIO_2_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:15]
  assign io_SRAMIO_3_cen = ~_T_4413; // @[Cache.scala 147:13]
  assign io_SRAMIO_3_wen = ~_T_4413; // @[Cache.scala 149:13]
  assign io_SRAMIO_3_wdata = io_cacheOut_r_last_i ? _T_4365 : _T_4366; // @[Cache.scala 150:15]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 148:14]
  assign io_SRAMIO_3_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cacheState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  vArrayWire_63_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vArrayWire_62_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  vArrayWire_61_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  vArrayWire_60_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vArrayWire_59_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  vArrayWire_58_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  vArrayWire_57_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  vArrayWire_56_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  vArrayWire_55_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  vArrayWire_54_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vArrayWire_53_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  vArrayWire_52_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  vArrayWire_51_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  vArrayWire_50_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  vArrayWire_49_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  vArrayWire_48_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  vArrayWire_47_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  vArrayWire_46_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  vArrayWire_45_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  vArrayWire_44_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  vArrayWire_43_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  vArrayWire_42_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  vArrayWire_41_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  vArrayWire_40_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  vArrayWire_39_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  vArrayWire_38_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vArrayWire_37_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  vArrayWire_36_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  vArrayWire_35_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  vArrayWire_34_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  vArrayWire_33_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  vArrayWire_32_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  vArrayWire_31_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  vArrayWire_30_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  vArrayWire_29_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  vArrayWire_28_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  vArrayWire_27_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  vArrayWire_26_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  vArrayWire_25_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  vArrayWire_24_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  vArrayWire_23_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  vArrayWire_22_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  vArrayWire_21_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  vArrayWire_20_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  vArrayWire_19_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  vArrayWire_18_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  vArrayWire_17_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  vArrayWire_16_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  vArrayWire_15_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  vArrayWire_14_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  vArrayWire_13_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  vArrayWire_12_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vArrayWire_11_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  vArrayWire_10_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  vArrayWire_9_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  vArrayWire_8_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  vArrayWire_7_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  vArrayWire_6_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  vArrayWire_5_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  vArrayWire_4_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  vArrayWire_3_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  vArrayWire_2_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  vArrayWire_1_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  vArrayWire_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tagArrayWire_63_0 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tagArrayWire_62_0 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tagArrayWire_61_0 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tagArrayWire_60_0 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tagArrayWire_59_0 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tagArrayWire_58_0 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tagArrayWire_57_0 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tagArrayWire_56_0 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tagArrayWire_55_0 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tagArrayWire_54_0 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tagArrayWire_53_0 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tagArrayWire_52_0 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tagArrayWire_51_0 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tagArrayWire_50_0 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tagArrayWire_49_0 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tagArrayWire_48_0 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tagArrayWire_47_0 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tagArrayWire_46_0 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tagArrayWire_45_0 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tagArrayWire_44_0 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tagArrayWire_43_0 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tagArrayWire_42_0 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tagArrayWire_41_0 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tagArrayWire_40_0 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tagArrayWire_39_0 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tagArrayWire_38_0 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tagArrayWire_37_0 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tagArrayWire_36_0 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tagArrayWire_35_0 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tagArrayWire_34_0 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tagArrayWire_33_0 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tagArrayWire_32_0 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tagArrayWire_31_0 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tagArrayWire_30_0 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tagArrayWire_29_0 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tagArrayWire_28_0 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tagArrayWire_27_0 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tagArrayWire_26_0 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tagArrayWire_25_0 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tagArrayWire_24_0 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tagArrayWire_23_0 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tagArrayWire_22_0 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tagArrayWire_21_0 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tagArrayWire_20_0 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tagArrayWire_19_0 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tagArrayWire_18_0 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tagArrayWire_17_0 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tagArrayWire_16_0 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tagArrayWire_15_0 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tagArrayWire_14_0 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tagArrayWire_13_0 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tagArrayWire_12_0 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tagArrayWire_11_0 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tagArrayWire_10_0 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tagArrayWire_9_0 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tagArrayWire_8_0 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tagArrayWire_7_0 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tagArrayWire_6_0 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tagArrayWire_5_0 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tagArrayWire_4_0 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tagArrayWire_3_0 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tagArrayWire_2_0 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tagArrayWire_1_0 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  tagArrayWire_0_0 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  vArrayWire_63_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  vArrayWire_62_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  vArrayWire_61_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  vArrayWire_60_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  vArrayWire_59_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  vArrayWire_58_1 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  vArrayWire_57_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  vArrayWire_56_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  vArrayWire_55_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  vArrayWire_54_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  vArrayWire_53_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  vArrayWire_52_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  vArrayWire_51_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  vArrayWire_50_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  vArrayWire_49_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  vArrayWire_48_1 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  vArrayWire_47_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  vArrayWire_46_1 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  vArrayWire_45_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  vArrayWire_44_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  vArrayWire_43_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  vArrayWire_42_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  vArrayWire_41_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  vArrayWire_40_1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  vArrayWire_39_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  vArrayWire_38_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  vArrayWire_37_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  vArrayWire_36_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  vArrayWire_35_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  vArrayWire_34_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  vArrayWire_33_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  vArrayWire_32_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  vArrayWire_31_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  vArrayWire_30_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  vArrayWire_29_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  vArrayWire_28_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  vArrayWire_27_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  vArrayWire_26_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  vArrayWire_25_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  vArrayWire_24_1 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  vArrayWire_23_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  vArrayWire_22_1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  vArrayWire_21_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  vArrayWire_20_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  vArrayWire_19_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  vArrayWire_18_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  vArrayWire_17_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  vArrayWire_16_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  vArrayWire_15_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  vArrayWire_14_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  vArrayWire_13_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  vArrayWire_12_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  vArrayWire_11_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  vArrayWire_10_1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vArrayWire_9_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  vArrayWire_8_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  vArrayWire_7_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  vArrayWire_6_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  vArrayWire_5_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  vArrayWire_4_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  vArrayWire_3_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  vArrayWire_2_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  vArrayWire_1_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  vArrayWire_0_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tagArrayWire_63_1 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  tagArrayWire_62_1 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  tagArrayWire_61_1 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  tagArrayWire_60_1 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  tagArrayWire_59_1 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  tagArrayWire_58_1 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  tagArrayWire_57_1 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  tagArrayWire_56_1 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  tagArrayWire_55_1 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  tagArrayWire_54_1 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  tagArrayWire_53_1 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  tagArrayWire_52_1 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  tagArrayWire_51_1 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  tagArrayWire_50_1 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  tagArrayWire_49_1 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  tagArrayWire_48_1 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  tagArrayWire_47_1 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  tagArrayWire_46_1 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  tagArrayWire_45_1 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  tagArrayWire_44_1 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  tagArrayWire_43_1 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  tagArrayWire_42_1 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  tagArrayWire_41_1 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  tagArrayWire_40_1 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  tagArrayWire_39_1 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  tagArrayWire_38_1 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  tagArrayWire_37_1 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  tagArrayWire_36_1 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  tagArrayWire_35_1 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  tagArrayWire_34_1 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  tagArrayWire_33_1 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  tagArrayWire_32_1 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  tagArrayWire_31_1 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  tagArrayWire_30_1 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  tagArrayWire_29_1 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  tagArrayWire_28_1 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  tagArrayWire_27_1 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  tagArrayWire_26_1 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  tagArrayWire_25_1 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  tagArrayWire_24_1 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  tagArrayWire_23_1 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  tagArrayWire_22_1 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  tagArrayWire_21_1 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  tagArrayWire_20_1 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  tagArrayWire_19_1 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  tagArrayWire_18_1 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  tagArrayWire_17_1 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  tagArrayWire_16_1 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  tagArrayWire_15_1 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  tagArrayWire_14_1 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  tagArrayWire_13_1 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  tagArrayWire_12_1 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  tagArrayWire_11_1 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  tagArrayWire_10_1 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  tagArrayWire_9_1 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  tagArrayWire_8_1 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  tagArrayWire_7_1 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  tagArrayWire_6_1 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  tagArrayWire_5_1 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  tagArrayWire_4_1 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  tagArrayWire_3_1 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  tagArrayWire_2_1 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  tagArrayWire_1_1 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  tagArrayWire_0_1 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  vArrayWire_63_2 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  vArrayWire_62_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  vArrayWire_61_2 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  vArrayWire_60_2 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  vArrayWire_59_2 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  vArrayWire_58_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  vArrayWire_57_2 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  vArrayWire_56_2 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  vArrayWire_55_2 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  vArrayWire_54_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  vArrayWire_53_2 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  vArrayWire_52_2 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  vArrayWire_51_2 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  vArrayWire_50_2 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  vArrayWire_49_2 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  vArrayWire_48_2 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  vArrayWire_47_2 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  vArrayWire_46_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  vArrayWire_45_2 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  vArrayWire_44_2 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  vArrayWire_43_2 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  vArrayWire_42_2 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  vArrayWire_41_2 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  vArrayWire_40_2 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  vArrayWire_39_2 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  vArrayWire_38_2 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  vArrayWire_37_2 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  vArrayWire_36_2 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  vArrayWire_35_2 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  vArrayWire_34_2 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  vArrayWire_33_2 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  vArrayWire_32_2 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  vArrayWire_31_2 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  vArrayWire_30_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  vArrayWire_29_2 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  vArrayWire_28_2 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  vArrayWire_27_2 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  vArrayWire_26_2 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  vArrayWire_25_2 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  vArrayWire_24_2 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  vArrayWire_23_2 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  vArrayWire_22_2 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  vArrayWire_21_2 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  vArrayWire_20_2 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  vArrayWire_19_2 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  vArrayWire_18_2 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  vArrayWire_17_2 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  vArrayWire_16_2 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  vArrayWire_15_2 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  vArrayWire_14_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  vArrayWire_13_2 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  vArrayWire_12_2 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  vArrayWire_11_2 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  vArrayWire_10_2 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  vArrayWire_9_2 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  vArrayWire_8_2 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  vArrayWire_7_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  vArrayWire_6_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  vArrayWire_5_2 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  vArrayWire_4_2 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  vArrayWire_3_2 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  vArrayWire_2_2 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  vArrayWire_1_2 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  vArrayWire_0_2 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  tagArrayWire_63_2 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  tagArrayWire_62_2 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  tagArrayWire_61_2 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  tagArrayWire_60_2 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  tagArrayWire_59_2 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  tagArrayWire_58_2 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  tagArrayWire_57_2 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  tagArrayWire_56_2 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  tagArrayWire_55_2 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  tagArrayWire_54_2 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  tagArrayWire_53_2 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  tagArrayWire_52_2 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  tagArrayWire_51_2 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  tagArrayWire_50_2 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  tagArrayWire_49_2 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  tagArrayWire_48_2 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  tagArrayWire_47_2 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  tagArrayWire_46_2 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  tagArrayWire_45_2 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  tagArrayWire_44_2 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  tagArrayWire_43_2 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  tagArrayWire_42_2 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  tagArrayWire_41_2 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  tagArrayWire_40_2 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  tagArrayWire_39_2 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  tagArrayWire_38_2 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  tagArrayWire_37_2 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  tagArrayWire_36_2 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  tagArrayWire_35_2 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  tagArrayWire_34_2 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  tagArrayWire_33_2 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  tagArrayWire_32_2 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  tagArrayWire_31_2 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  tagArrayWire_30_2 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  tagArrayWire_29_2 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  tagArrayWire_28_2 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  tagArrayWire_27_2 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  tagArrayWire_26_2 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  tagArrayWire_25_2 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  tagArrayWire_24_2 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  tagArrayWire_23_2 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  tagArrayWire_22_2 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  tagArrayWire_21_2 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  tagArrayWire_20_2 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  tagArrayWire_19_2 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  tagArrayWire_18_2 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  tagArrayWire_17_2 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  tagArrayWire_16_2 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  tagArrayWire_15_2 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  tagArrayWire_14_2 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  tagArrayWire_13_2 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  tagArrayWire_12_2 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  tagArrayWire_11_2 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  tagArrayWire_10_2 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  tagArrayWire_9_2 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  tagArrayWire_8_2 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  tagArrayWire_7_2 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  tagArrayWire_6_2 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  tagArrayWire_5_2 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  tagArrayWire_4_2 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  tagArrayWire_3_2 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  tagArrayWire_2_2 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  tagArrayWire_1_2 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  tagArrayWire_0_2 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  vArrayWire_63_3 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  vArrayWire_62_3 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  vArrayWire_61_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  vArrayWire_60_3 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  vArrayWire_59_3 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  vArrayWire_58_3 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  vArrayWire_57_3 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  vArrayWire_56_3 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  vArrayWire_55_3 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  vArrayWire_54_3 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  vArrayWire_53_3 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  vArrayWire_52_3 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  vArrayWire_51_3 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  vArrayWire_50_3 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  vArrayWire_49_3 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  vArrayWire_48_3 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  vArrayWire_47_3 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  vArrayWire_46_3 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  vArrayWire_45_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  vArrayWire_44_3 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  vArrayWire_43_3 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  vArrayWire_42_3 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  vArrayWire_41_3 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  vArrayWire_40_3 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  vArrayWire_39_3 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  vArrayWire_38_3 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  vArrayWire_37_3 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  vArrayWire_36_3 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  vArrayWire_35_3 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  vArrayWire_34_3 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  vArrayWire_33_3 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  vArrayWire_32_3 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  vArrayWire_31_3 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  vArrayWire_30_3 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  vArrayWire_29_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  vArrayWire_28_3 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  vArrayWire_27_3 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  vArrayWire_26_3 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  vArrayWire_25_3 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  vArrayWire_24_3 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  vArrayWire_23_3 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  vArrayWire_22_3 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  vArrayWire_21_3 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  vArrayWire_20_3 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  vArrayWire_19_3 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  vArrayWire_18_3 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  vArrayWire_17_3 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  vArrayWire_16_3 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  vArrayWire_15_3 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  vArrayWire_14_3 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  vArrayWire_13_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  vArrayWire_12_3 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  vArrayWire_11_3 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  vArrayWire_10_3 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  vArrayWire_9_3 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  vArrayWire_8_3 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  vArrayWire_7_3 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  vArrayWire_6_3 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  vArrayWire_5_3 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  vArrayWire_4_3 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  vArrayWire_3_3 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  vArrayWire_2_3 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  vArrayWire_1_3 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  vArrayWire_0_3 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  tagArrayWire_63_3 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  tagArrayWire_62_3 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  tagArrayWire_61_3 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  tagArrayWire_60_3 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  tagArrayWire_59_3 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  tagArrayWire_58_3 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  tagArrayWire_57_3 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  tagArrayWire_56_3 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  tagArrayWire_55_3 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  tagArrayWire_54_3 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  tagArrayWire_53_3 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  tagArrayWire_52_3 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  tagArrayWire_51_3 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  tagArrayWire_50_3 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  tagArrayWire_49_3 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  tagArrayWire_48_3 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  tagArrayWire_47_3 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  tagArrayWire_46_3 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  tagArrayWire_45_3 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  tagArrayWire_44_3 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  tagArrayWire_43_3 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  tagArrayWire_42_3 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  tagArrayWire_41_3 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  tagArrayWire_40_3 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  tagArrayWire_39_3 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  tagArrayWire_38_3 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  tagArrayWire_37_3 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  tagArrayWire_36_3 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  tagArrayWire_35_3 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  tagArrayWire_34_3 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  tagArrayWire_33_3 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  tagArrayWire_32_3 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  tagArrayWire_31_3 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  tagArrayWire_30_3 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  tagArrayWire_29_3 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  tagArrayWire_28_3 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  tagArrayWire_27_3 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  tagArrayWire_26_3 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  tagArrayWire_25_3 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  tagArrayWire_24_3 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  tagArrayWire_23_3 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  tagArrayWire_22_3 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  tagArrayWire_21_3 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  tagArrayWire_20_3 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  tagArrayWire_19_3 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  tagArrayWire_18_3 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  tagArrayWire_17_3 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  tagArrayWire_16_3 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  tagArrayWire_15_3 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  tagArrayWire_14_3 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  tagArrayWire_13_3 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  tagArrayWire_12_3 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  tagArrayWire_11_3 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  tagArrayWire_10_3 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  tagArrayWire_9_3 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  tagArrayWire_8_3 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  tagArrayWire_7_3 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  tagArrayWire_6_3 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  tagArrayWire_5_3 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  tagArrayWire_4_3 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  tagArrayWire_3_3 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  tagArrayWire_2_3 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  tagArrayWire_1_3 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  tagArrayWire_0_3 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  selArrayWire_1 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  selArrayWire_0 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  selArrayWire_2 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  selArrayWire_3 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  selArrayWire_4 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  selArrayWire_5 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  selArrayWire_6 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  selArrayWire_7 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  selArrayWire_8 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  selArrayWire_9 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  selArrayWire_10 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  selArrayWire_11 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  selArrayWire_12 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  selArrayWire_13 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  selArrayWire_14 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  selArrayWire_15 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  selArrayWire_16 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  selArrayWire_17 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  selArrayWire_18 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  selArrayWire_19 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  selArrayWire_20 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  selArrayWire_21 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  selArrayWire_22 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  selArrayWire_23 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  selArrayWire_24 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  selArrayWire_25 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  selArrayWire_26 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  selArrayWire_27 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  selArrayWire_28 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  selArrayWire_29 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  selArrayWire_30 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  selArrayWire_31 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  selArrayWire_32 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  selArrayWire_33 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  selArrayWire_34 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  selArrayWire_35 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  selArrayWire_36 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  selArrayWire_37 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  selArrayWire_38 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  selArrayWire_39 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  selArrayWire_40 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  selArrayWire_41 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  selArrayWire_42 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  selArrayWire_43 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  selArrayWire_44 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  selArrayWire_45 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  selArrayWire_46 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  selArrayWire_47 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  selArrayWire_48 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  selArrayWire_49 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  selArrayWire_50 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  selArrayWire_51 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  selArrayWire_52 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  selArrayWire_53 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  selArrayWire_54 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  selArrayWire_55 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  selArrayWire_56 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  selArrayWire_57 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  selArrayWire_58 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  selArrayWire_59 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  selArrayWire_60 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  selArrayWire_61 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  selArrayWire_62 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  selArrayWire_63 = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cacheState <= 1'h0;
    end else if (cacheState) begin
      if (io_cacheOut_r_last_i) begin
        cacheState <= 1'h0;
      end else begin
        cacheState <= 1'h1;
      end
    end else begin
      cacheState <= IdleMux;
    end
    if (_T_412) begin
      vArrayWire_63_0 <= 1'h0;
    end else begin
      vArrayWire_63_0 <= _GEN_569;
    end
    if (_T_412) begin
      vArrayWire_62_0 <= 1'h0;
    end else begin
      vArrayWire_62_0 <= _GEN_560;
    end
    if (_T_412) begin
      vArrayWire_61_0 <= 1'h0;
    end else begin
      vArrayWire_61_0 <= _GEN_551;
    end
    if (_T_412) begin
      vArrayWire_60_0 <= 1'h0;
    end else begin
      vArrayWire_60_0 <= _GEN_542;
    end
    if (_T_412) begin
      vArrayWire_59_0 <= 1'h0;
    end else begin
      vArrayWire_59_0 <= _GEN_533;
    end
    if (_T_412) begin
      vArrayWire_58_0 <= 1'h0;
    end else begin
      vArrayWire_58_0 <= _GEN_524;
    end
    if (_T_412) begin
      vArrayWire_57_0 <= 1'h0;
    end else begin
      vArrayWire_57_0 <= _GEN_515;
    end
    if (_T_412) begin
      vArrayWire_56_0 <= 1'h0;
    end else begin
      vArrayWire_56_0 <= _GEN_506;
    end
    if (_T_412) begin
      vArrayWire_55_0 <= 1'h0;
    end else begin
      vArrayWire_55_0 <= _GEN_497;
    end
    if (_T_412) begin
      vArrayWire_54_0 <= 1'h0;
    end else begin
      vArrayWire_54_0 <= _GEN_488;
    end
    if (_T_412) begin
      vArrayWire_53_0 <= 1'h0;
    end else begin
      vArrayWire_53_0 <= _GEN_479;
    end
    if (_T_412) begin
      vArrayWire_52_0 <= 1'h0;
    end else begin
      vArrayWire_52_0 <= _GEN_470;
    end
    if (_T_412) begin
      vArrayWire_51_0 <= 1'h0;
    end else begin
      vArrayWire_51_0 <= _GEN_461;
    end
    if (_T_412) begin
      vArrayWire_50_0 <= 1'h0;
    end else begin
      vArrayWire_50_0 <= _GEN_452;
    end
    if (_T_412) begin
      vArrayWire_49_0 <= 1'h0;
    end else begin
      vArrayWire_49_0 <= _GEN_443;
    end
    if (_T_412) begin
      vArrayWire_48_0 <= 1'h0;
    end else begin
      vArrayWire_48_0 <= _GEN_434;
    end
    if (_T_412) begin
      vArrayWire_47_0 <= 1'h0;
    end else begin
      vArrayWire_47_0 <= _GEN_425;
    end
    if (_T_412) begin
      vArrayWire_46_0 <= 1'h0;
    end else begin
      vArrayWire_46_0 <= _GEN_416;
    end
    if (_T_412) begin
      vArrayWire_45_0 <= 1'h0;
    end else begin
      vArrayWire_45_0 <= _GEN_407;
    end
    if (_T_412) begin
      vArrayWire_44_0 <= 1'h0;
    end else begin
      vArrayWire_44_0 <= _GEN_398;
    end
    if (_T_412) begin
      vArrayWire_43_0 <= 1'h0;
    end else begin
      vArrayWire_43_0 <= _GEN_389;
    end
    if (_T_412) begin
      vArrayWire_42_0 <= 1'h0;
    end else begin
      vArrayWire_42_0 <= _GEN_380;
    end
    if (_T_412) begin
      vArrayWire_41_0 <= 1'h0;
    end else begin
      vArrayWire_41_0 <= _GEN_371;
    end
    if (_T_412) begin
      vArrayWire_40_0 <= 1'h0;
    end else begin
      vArrayWire_40_0 <= _GEN_362;
    end
    if (_T_412) begin
      vArrayWire_39_0 <= 1'h0;
    end else begin
      vArrayWire_39_0 <= _GEN_353;
    end
    if (_T_412) begin
      vArrayWire_38_0 <= 1'h0;
    end else begin
      vArrayWire_38_0 <= _GEN_344;
    end
    if (_T_412) begin
      vArrayWire_37_0 <= 1'h0;
    end else begin
      vArrayWire_37_0 <= _GEN_335;
    end
    if (_T_412) begin
      vArrayWire_36_0 <= 1'h0;
    end else begin
      vArrayWire_36_0 <= _GEN_326;
    end
    if (_T_412) begin
      vArrayWire_35_0 <= 1'h0;
    end else begin
      vArrayWire_35_0 <= _GEN_317;
    end
    if (_T_412) begin
      vArrayWire_34_0 <= 1'h0;
    end else begin
      vArrayWire_34_0 <= _GEN_308;
    end
    if (_T_412) begin
      vArrayWire_33_0 <= 1'h0;
    end else begin
      vArrayWire_33_0 <= _GEN_299;
    end
    if (_T_412) begin
      vArrayWire_32_0 <= 1'h0;
    end else begin
      vArrayWire_32_0 <= _GEN_290;
    end
    if (_T_412) begin
      vArrayWire_31_0 <= 1'h0;
    end else begin
      vArrayWire_31_0 <= _GEN_281;
    end
    if (_T_412) begin
      vArrayWire_30_0 <= 1'h0;
    end else begin
      vArrayWire_30_0 <= _GEN_272;
    end
    if (_T_412) begin
      vArrayWire_29_0 <= 1'h0;
    end else begin
      vArrayWire_29_0 <= _GEN_263;
    end
    if (_T_412) begin
      vArrayWire_28_0 <= 1'h0;
    end else begin
      vArrayWire_28_0 <= _GEN_254;
    end
    if (_T_412) begin
      vArrayWire_27_0 <= 1'h0;
    end else begin
      vArrayWire_27_0 <= _GEN_245;
    end
    if (_T_412) begin
      vArrayWire_26_0 <= 1'h0;
    end else begin
      vArrayWire_26_0 <= _GEN_236;
    end
    if (_T_412) begin
      vArrayWire_25_0 <= 1'h0;
    end else begin
      vArrayWire_25_0 <= _GEN_227;
    end
    if (_T_412) begin
      vArrayWire_24_0 <= 1'h0;
    end else begin
      vArrayWire_24_0 <= _GEN_218;
    end
    if (_T_412) begin
      vArrayWire_23_0 <= 1'h0;
    end else begin
      vArrayWire_23_0 <= _GEN_209;
    end
    if (_T_412) begin
      vArrayWire_22_0 <= 1'h0;
    end else begin
      vArrayWire_22_0 <= _GEN_200;
    end
    if (_T_412) begin
      vArrayWire_21_0 <= 1'h0;
    end else begin
      vArrayWire_21_0 <= _GEN_191;
    end
    if (_T_412) begin
      vArrayWire_20_0 <= 1'h0;
    end else begin
      vArrayWire_20_0 <= _GEN_182;
    end
    if (_T_412) begin
      vArrayWire_19_0 <= 1'h0;
    end else begin
      vArrayWire_19_0 <= _GEN_173;
    end
    if (_T_412) begin
      vArrayWire_18_0 <= 1'h0;
    end else begin
      vArrayWire_18_0 <= _GEN_164;
    end
    if (_T_412) begin
      vArrayWire_17_0 <= 1'h0;
    end else begin
      vArrayWire_17_0 <= _GEN_155;
    end
    if (_T_412) begin
      vArrayWire_16_0 <= 1'h0;
    end else begin
      vArrayWire_16_0 <= _GEN_146;
    end
    if (_T_412) begin
      vArrayWire_15_0 <= 1'h0;
    end else begin
      vArrayWire_15_0 <= _GEN_137;
    end
    if (_T_412) begin
      vArrayWire_14_0 <= 1'h0;
    end else begin
      vArrayWire_14_0 <= _GEN_128;
    end
    if (_T_412) begin
      vArrayWire_13_0 <= 1'h0;
    end else begin
      vArrayWire_13_0 <= _GEN_119;
    end
    if (_T_412) begin
      vArrayWire_12_0 <= 1'h0;
    end else begin
      vArrayWire_12_0 <= _GEN_110;
    end
    if (_T_412) begin
      vArrayWire_11_0 <= 1'h0;
    end else begin
      vArrayWire_11_0 <= _GEN_101;
    end
    if (_T_412) begin
      vArrayWire_10_0 <= 1'h0;
    end else begin
      vArrayWire_10_0 <= _GEN_92;
    end
    if (_T_412) begin
      vArrayWire_9_0 <= 1'h0;
    end else begin
      vArrayWire_9_0 <= _GEN_83;
    end
    if (_T_412) begin
      vArrayWire_8_0 <= 1'h0;
    end else begin
      vArrayWire_8_0 <= _GEN_74;
    end
    if (_T_412) begin
      vArrayWire_7_0 <= 1'h0;
    end else begin
      vArrayWire_7_0 <= _GEN_65;
    end
    if (_T_412) begin
      vArrayWire_6_0 <= 1'h0;
    end else begin
      vArrayWire_6_0 <= _GEN_56;
    end
    if (_T_412) begin
      vArrayWire_5_0 <= 1'h0;
    end else begin
      vArrayWire_5_0 <= _GEN_47;
    end
    if (_T_412) begin
      vArrayWire_4_0 <= 1'h0;
    end else begin
      vArrayWire_4_0 <= _GEN_38;
    end
    if (_T_412) begin
      vArrayWire_3_0 <= 1'h0;
    end else begin
      vArrayWire_3_0 <= _GEN_29;
    end
    if (_T_412) begin
      vArrayWire_2_0 <= 1'h0;
    end else begin
      vArrayWire_2_0 <= _GEN_20;
    end
    if (_T_412) begin
      vArrayWire_1_0 <= 1'h0;
    end else begin
      vArrayWire_1_0 <= _GEN_11;
    end
    if (_T_412) begin
      vArrayWire_0_0 <= 1'h0;
    end else begin
      vArrayWire_0_0 <= _GEN_2;
    end
    if (reset) begin
      tagArrayWire_63_0 <= 22'h0;
    end else if (_T_4252) begin
      tagArrayWire_63_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_0 <= 22'h0;
    end else if (_T_4191) begin
      tagArrayWire_62_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_0 <= 22'h0;
    end else if (_T_4130) begin
      tagArrayWire_61_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_0 <= 22'h0;
    end else if (_T_4069) begin
      tagArrayWire_60_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_0 <= 22'h0;
    end else if (_T_4008) begin
      tagArrayWire_59_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_0 <= 22'h0;
    end else if (_T_3947) begin
      tagArrayWire_58_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_0 <= 22'h0;
    end else if (_T_3886) begin
      tagArrayWire_57_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_0 <= 22'h0;
    end else if (_T_3825) begin
      tagArrayWire_56_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_0 <= 22'h0;
    end else if (_T_3764) begin
      tagArrayWire_55_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_0 <= 22'h0;
    end else if (_T_3703) begin
      tagArrayWire_54_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_0 <= 22'h0;
    end else if (_T_3642) begin
      tagArrayWire_53_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_0 <= 22'h0;
    end else if (_T_3581) begin
      tagArrayWire_52_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_0 <= 22'h0;
    end else if (_T_3520) begin
      tagArrayWire_51_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_0 <= 22'h0;
    end else if (_T_3459) begin
      tagArrayWire_50_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_0 <= 22'h0;
    end else if (_T_3398) begin
      tagArrayWire_49_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_0 <= 22'h0;
    end else if (_T_3337) begin
      tagArrayWire_48_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_0 <= 22'h0;
    end else if (_T_3276) begin
      tagArrayWire_47_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_0 <= 22'h0;
    end else if (_T_3215) begin
      tagArrayWire_46_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_0 <= 22'h0;
    end else if (_T_3154) begin
      tagArrayWire_45_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_0 <= 22'h0;
    end else if (_T_3093) begin
      tagArrayWire_44_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_0 <= 22'h0;
    end else if (_T_3032) begin
      tagArrayWire_43_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_0 <= 22'h0;
    end else if (_T_2971) begin
      tagArrayWire_42_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_0 <= 22'h0;
    end else if (_T_2910) begin
      tagArrayWire_41_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_0 <= 22'h0;
    end else if (_T_2849) begin
      tagArrayWire_40_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_0 <= 22'h0;
    end else if (_T_2788) begin
      tagArrayWire_39_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_0 <= 22'h0;
    end else if (_T_2727) begin
      tagArrayWire_38_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_0 <= 22'h0;
    end else if (_T_2666) begin
      tagArrayWire_37_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_0 <= 22'h0;
    end else if (_T_2605) begin
      tagArrayWire_36_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_0 <= 22'h0;
    end else if (_T_2544) begin
      tagArrayWire_35_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_0 <= 22'h0;
    end else if (_T_2483) begin
      tagArrayWire_34_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_0 <= 22'h0;
    end else if (_T_2422) begin
      tagArrayWire_33_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_0 <= 22'h0;
    end else if (_T_2361) begin
      tagArrayWire_32_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_0 <= 22'h0;
    end else if (_T_2300) begin
      tagArrayWire_31_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_0 <= 22'h0;
    end else if (_T_2239) begin
      tagArrayWire_30_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_0 <= 22'h0;
    end else if (_T_2178) begin
      tagArrayWire_29_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_0 <= 22'h0;
    end else if (_T_2117) begin
      tagArrayWire_28_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_0 <= 22'h0;
    end else if (_T_2056) begin
      tagArrayWire_27_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_0 <= 22'h0;
    end else if (_T_1995) begin
      tagArrayWire_26_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_0 <= 22'h0;
    end else if (_T_1934) begin
      tagArrayWire_25_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_0 <= 22'h0;
    end else if (_T_1873) begin
      tagArrayWire_24_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_0 <= 22'h0;
    end else if (_T_1812) begin
      tagArrayWire_23_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_0 <= 22'h0;
    end else if (_T_1751) begin
      tagArrayWire_22_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_0 <= 22'h0;
    end else if (_T_1690) begin
      tagArrayWire_21_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_0 <= 22'h0;
    end else if (_T_1629) begin
      tagArrayWire_20_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_0 <= 22'h0;
    end else if (_T_1568) begin
      tagArrayWire_19_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_0 <= 22'h0;
    end else if (_T_1507) begin
      tagArrayWire_18_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_0 <= 22'h0;
    end else if (_T_1446) begin
      tagArrayWire_17_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_0 <= 22'h0;
    end else if (_T_1385) begin
      tagArrayWire_16_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_0 <= 22'h0;
    end else if (_T_1324) begin
      tagArrayWire_15_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_0 <= 22'h0;
    end else if (_T_1263) begin
      tagArrayWire_14_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_0 <= 22'h0;
    end else if (_T_1202) begin
      tagArrayWire_13_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_0 <= 22'h0;
    end else if (_T_1141) begin
      tagArrayWire_12_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_0 <= 22'h0;
    end else if (_T_1080) begin
      tagArrayWire_11_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_0 <= 22'h0;
    end else if (_T_1019) begin
      tagArrayWire_10_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_0 <= 22'h0;
    end else if (_T_958) begin
      tagArrayWire_9_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_0 <= 22'h0;
    end else if (_T_897) begin
      tagArrayWire_8_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_0 <= 22'h0;
    end else if (_T_836) begin
      tagArrayWire_7_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_0 <= 22'h0;
    end else if (_T_775) begin
      tagArrayWire_6_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_0 <= 22'h0;
    end else if (_T_714) begin
      tagArrayWire_5_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_0 <= 22'h0;
    end else if (_T_653) begin
      tagArrayWire_4_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_0 <= 22'h0;
    end else if (_T_592) begin
      tagArrayWire_3_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_0 <= 22'h0;
    end else if (_T_531) begin
      tagArrayWire_2_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_0 <= 22'h0;
    end else if (_T_470) begin
      tagArrayWire_1_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_0 <= 22'h0;
    end else if (_T_409) begin
      tagArrayWire_0_0 <= tag;
    end
    if (_T_412) begin
      vArrayWire_63_1 <= 1'h0;
    end else begin
      vArrayWire_63_1 <= _GEN_571;
    end
    if (_T_412) begin
      vArrayWire_62_1 <= 1'h0;
    end else begin
      vArrayWire_62_1 <= _GEN_562;
    end
    if (_T_412) begin
      vArrayWire_61_1 <= 1'h0;
    end else begin
      vArrayWire_61_1 <= _GEN_553;
    end
    if (_T_412) begin
      vArrayWire_60_1 <= 1'h0;
    end else begin
      vArrayWire_60_1 <= _GEN_544;
    end
    if (_T_412) begin
      vArrayWire_59_1 <= 1'h0;
    end else begin
      vArrayWire_59_1 <= _GEN_535;
    end
    if (_T_412) begin
      vArrayWire_58_1 <= 1'h0;
    end else begin
      vArrayWire_58_1 <= _GEN_526;
    end
    if (_T_412) begin
      vArrayWire_57_1 <= 1'h0;
    end else begin
      vArrayWire_57_1 <= _GEN_517;
    end
    if (_T_412) begin
      vArrayWire_56_1 <= 1'h0;
    end else begin
      vArrayWire_56_1 <= _GEN_508;
    end
    if (_T_412) begin
      vArrayWire_55_1 <= 1'h0;
    end else begin
      vArrayWire_55_1 <= _GEN_499;
    end
    if (_T_412) begin
      vArrayWire_54_1 <= 1'h0;
    end else begin
      vArrayWire_54_1 <= _GEN_490;
    end
    if (_T_412) begin
      vArrayWire_53_1 <= 1'h0;
    end else begin
      vArrayWire_53_1 <= _GEN_481;
    end
    if (_T_412) begin
      vArrayWire_52_1 <= 1'h0;
    end else begin
      vArrayWire_52_1 <= _GEN_472;
    end
    if (_T_412) begin
      vArrayWire_51_1 <= 1'h0;
    end else begin
      vArrayWire_51_1 <= _GEN_463;
    end
    if (_T_412) begin
      vArrayWire_50_1 <= 1'h0;
    end else begin
      vArrayWire_50_1 <= _GEN_454;
    end
    if (_T_412) begin
      vArrayWire_49_1 <= 1'h0;
    end else begin
      vArrayWire_49_1 <= _GEN_445;
    end
    if (_T_412) begin
      vArrayWire_48_1 <= 1'h0;
    end else begin
      vArrayWire_48_1 <= _GEN_436;
    end
    if (_T_412) begin
      vArrayWire_47_1 <= 1'h0;
    end else begin
      vArrayWire_47_1 <= _GEN_427;
    end
    if (_T_412) begin
      vArrayWire_46_1 <= 1'h0;
    end else begin
      vArrayWire_46_1 <= _GEN_418;
    end
    if (_T_412) begin
      vArrayWire_45_1 <= 1'h0;
    end else begin
      vArrayWire_45_1 <= _GEN_409;
    end
    if (_T_412) begin
      vArrayWire_44_1 <= 1'h0;
    end else begin
      vArrayWire_44_1 <= _GEN_400;
    end
    if (_T_412) begin
      vArrayWire_43_1 <= 1'h0;
    end else begin
      vArrayWire_43_1 <= _GEN_391;
    end
    if (_T_412) begin
      vArrayWire_42_1 <= 1'h0;
    end else begin
      vArrayWire_42_1 <= _GEN_382;
    end
    if (_T_412) begin
      vArrayWire_41_1 <= 1'h0;
    end else begin
      vArrayWire_41_1 <= _GEN_373;
    end
    if (_T_412) begin
      vArrayWire_40_1 <= 1'h0;
    end else begin
      vArrayWire_40_1 <= _GEN_364;
    end
    if (_T_412) begin
      vArrayWire_39_1 <= 1'h0;
    end else begin
      vArrayWire_39_1 <= _GEN_355;
    end
    if (_T_412) begin
      vArrayWire_38_1 <= 1'h0;
    end else begin
      vArrayWire_38_1 <= _GEN_346;
    end
    if (_T_412) begin
      vArrayWire_37_1 <= 1'h0;
    end else begin
      vArrayWire_37_1 <= _GEN_337;
    end
    if (_T_412) begin
      vArrayWire_36_1 <= 1'h0;
    end else begin
      vArrayWire_36_1 <= _GEN_328;
    end
    if (_T_412) begin
      vArrayWire_35_1 <= 1'h0;
    end else begin
      vArrayWire_35_1 <= _GEN_319;
    end
    if (_T_412) begin
      vArrayWire_34_1 <= 1'h0;
    end else begin
      vArrayWire_34_1 <= _GEN_310;
    end
    if (_T_412) begin
      vArrayWire_33_1 <= 1'h0;
    end else begin
      vArrayWire_33_1 <= _GEN_301;
    end
    if (_T_412) begin
      vArrayWire_32_1 <= 1'h0;
    end else begin
      vArrayWire_32_1 <= _GEN_292;
    end
    if (_T_412) begin
      vArrayWire_31_1 <= 1'h0;
    end else begin
      vArrayWire_31_1 <= _GEN_283;
    end
    if (_T_412) begin
      vArrayWire_30_1 <= 1'h0;
    end else begin
      vArrayWire_30_1 <= _GEN_274;
    end
    if (_T_412) begin
      vArrayWire_29_1 <= 1'h0;
    end else begin
      vArrayWire_29_1 <= _GEN_265;
    end
    if (_T_412) begin
      vArrayWire_28_1 <= 1'h0;
    end else begin
      vArrayWire_28_1 <= _GEN_256;
    end
    if (_T_412) begin
      vArrayWire_27_1 <= 1'h0;
    end else begin
      vArrayWire_27_1 <= _GEN_247;
    end
    if (_T_412) begin
      vArrayWire_26_1 <= 1'h0;
    end else begin
      vArrayWire_26_1 <= _GEN_238;
    end
    if (_T_412) begin
      vArrayWire_25_1 <= 1'h0;
    end else begin
      vArrayWire_25_1 <= _GEN_229;
    end
    if (_T_412) begin
      vArrayWire_24_1 <= 1'h0;
    end else begin
      vArrayWire_24_1 <= _GEN_220;
    end
    if (_T_412) begin
      vArrayWire_23_1 <= 1'h0;
    end else begin
      vArrayWire_23_1 <= _GEN_211;
    end
    if (_T_412) begin
      vArrayWire_22_1 <= 1'h0;
    end else begin
      vArrayWire_22_1 <= _GEN_202;
    end
    if (_T_412) begin
      vArrayWire_21_1 <= 1'h0;
    end else begin
      vArrayWire_21_1 <= _GEN_193;
    end
    if (_T_412) begin
      vArrayWire_20_1 <= 1'h0;
    end else begin
      vArrayWire_20_1 <= _GEN_184;
    end
    if (_T_412) begin
      vArrayWire_19_1 <= 1'h0;
    end else begin
      vArrayWire_19_1 <= _GEN_175;
    end
    if (_T_412) begin
      vArrayWire_18_1 <= 1'h0;
    end else begin
      vArrayWire_18_1 <= _GEN_166;
    end
    if (_T_412) begin
      vArrayWire_17_1 <= 1'h0;
    end else begin
      vArrayWire_17_1 <= _GEN_157;
    end
    if (_T_412) begin
      vArrayWire_16_1 <= 1'h0;
    end else begin
      vArrayWire_16_1 <= _GEN_148;
    end
    if (_T_412) begin
      vArrayWire_15_1 <= 1'h0;
    end else begin
      vArrayWire_15_1 <= _GEN_139;
    end
    if (_T_412) begin
      vArrayWire_14_1 <= 1'h0;
    end else begin
      vArrayWire_14_1 <= _GEN_130;
    end
    if (_T_412) begin
      vArrayWire_13_1 <= 1'h0;
    end else begin
      vArrayWire_13_1 <= _GEN_121;
    end
    if (_T_412) begin
      vArrayWire_12_1 <= 1'h0;
    end else begin
      vArrayWire_12_1 <= _GEN_112;
    end
    if (_T_412) begin
      vArrayWire_11_1 <= 1'h0;
    end else begin
      vArrayWire_11_1 <= _GEN_103;
    end
    if (_T_412) begin
      vArrayWire_10_1 <= 1'h0;
    end else begin
      vArrayWire_10_1 <= _GEN_94;
    end
    if (_T_412) begin
      vArrayWire_9_1 <= 1'h0;
    end else begin
      vArrayWire_9_1 <= _GEN_85;
    end
    if (_T_412) begin
      vArrayWire_8_1 <= 1'h0;
    end else begin
      vArrayWire_8_1 <= _GEN_76;
    end
    if (_T_412) begin
      vArrayWire_7_1 <= 1'h0;
    end else begin
      vArrayWire_7_1 <= _GEN_67;
    end
    if (_T_412) begin
      vArrayWire_6_1 <= 1'h0;
    end else begin
      vArrayWire_6_1 <= _GEN_58;
    end
    if (_T_412) begin
      vArrayWire_5_1 <= 1'h0;
    end else begin
      vArrayWire_5_1 <= _GEN_49;
    end
    if (_T_412) begin
      vArrayWire_4_1 <= 1'h0;
    end else begin
      vArrayWire_4_1 <= _GEN_40;
    end
    if (_T_412) begin
      vArrayWire_3_1 <= 1'h0;
    end else begin
      vArrayWire_3_1 <= _GEN_31;
    end
    if (_T_412) begin
      vArrayWire_2_1 <= 1'h0;
    end else begin
      vArrayWire_2_1 <= _GEN_22;
    end
    if (_T_412) begin
      vArrayWire_1_1 <= 1'h0;
    end else begin
      vArrayWire_1_1 <= _GEN_13;
    end
    if (_T_412) begin
      vArrayWire_0_1 <= 1'h0;
    end else begin
      vArrayWire_0_1 <= _GEN_4;
    end
    if (reset) begin
      tagArrayWire_63_1 <= 22'h0;
    end else if (_T_4266) begin
      tagArrayWire_63_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_1 <= 22'h0;
    end else if (_T_4205) begin
      tagArrayWire_62_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_1 <= 22'h0;
    end else if (_T_4144) begin
      tagArrayWire_61_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_1 <= 22'h0;
    end else if (_T_4083) begin
      tagArrayWire_60_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_1 <= 22'h0;
    end else if (_T_4022) begin
      tagArrayWire_59_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_1 <= 22'h0;
    end else if (_T_3961) begin
      tagArrayWire_58_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_1 <= 22'h0;
    end else if (_T_3900) begin
      tagArrayWire_57_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_1 <= 22'h0;
    end else if (_T_3839) begin
      tagArrayWire_56_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_1 <= 22'h0;
    end else if (_T_3778) begin
      tagArrayWire_55_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_1 <= 22'h0;
    end else if (_T_3717) begin
      tagArrayWire_54_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_1 <= 22'h0;
    end else if (_T_3656) begin
      tagArrayWire_53_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_1 <= 22'h0;
    end else if (_T_3595) begin
      tagArrayWire_52_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_1 <= 22'h0;
    end else if (_T_3534) begin
      tagArrayWire_51_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_1 <= 22'h0;
    end else if (_T_3473) begin
      tagArrayWire_50_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_1 <= 22'h0;
    end else if (_T_3412) begin
      tagArrayWire_49_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_1 <= 22'h0;
    end else if (_T_3351) begin
      tagArrayWire_48_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_1 <= 22'h0;
    end else if (_T_3290) begin
      tagArrayWire_47_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_1 <= 22'h0;
    end else if (_T_3229) begin
      tagArrayWire_46_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_1 <= 22'h0;
    end else if (_T_3168) begin
      tagArrayWire_45_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_1 <= 22'h0;
    end else if (_T_3107) begin
      tagArrayWire_44_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_1 <= 22'h0;
    end else if (_T_3046) begin
      tagArrayWire_43_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_1 <= 22'h0;
    end else if (_T_2985) begin
      tagArrayWire_42_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_1 <= 22'h0;
    end else if (_T_2924) begin
      tagArrayWire_41_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_1 <= 22'h0;
    end else if (_T_2863) begin
      tagArrayWire_40_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_1 <= 22'h0;
    end else if (_T_2802) begin
      tagArrayWire_39_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_1 <= 22'h0;
    end else if (_T_2741) begin
      tagArrayWire_38_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_1 <= 22'h0;
    end else if (_T_2680) begin
      tagArrayWire_37_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_1 <= 22'h0;
    end else if (_T_2619) begin
      tagArrayWire_36_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_1 <= 22'h0;
    end else if (_T_2558) begin
      tagArrayWire_35_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_1 <= 22'h0;
    end else if (_T_2497) begin
      tagArrayWire_34_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_1 <= 22'h0;
    end else if (_T_2436) begin
      tagArrayWire_33_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_1 <= 22'h0;
    end else if (_T_2375) begin
      tagArrayWire_32_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_1 <= 22'h0;
    end else if (_T_2314) begin
      tagArrayWire_31_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_1 <= 22'h0;
    end else if (_T_2253) begin
      tagArrayWire_30_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_1 <= 22'h0;
    end else if (_T_2192) begin
      tagArrayWire_29_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_1 <= 22'h0;
    end else if (_T_2131) begin
      tagArrayWire_28_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_1 <= 22'h0;
    end else if (_T_2070) begin
      tagArrayWire_27_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_1 <= 22'h0;
    end else if (_T_2009) begin
      tagArrayWire_26_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_1 <= 22'h0;
    end else if (_T_1948) begin
      tagArrayWire_25_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_1 <= 22'h0;
    end else if (_T_1887) begin
      tagArrayWire_24_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_1 <= 22'h0;
    end else if (_T_1826) begin
      tagArrayWire_23_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_1 <= 22'h0;
    end else if (_T_1765) begin
      tagArrayWire_22_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_1 <= 22'h0;
    end else if (_T_1704) begin
      tagArrayWire_21_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_1 <= 22'h0;
    end else if (_T_1643) begin
      tagArrayWire_20_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_1 <= 22'h0;
    end else if (_T_1582) begin
      tagArrayWire_19_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_1 <= 22'h0;
    end else if (_T_1521) begin
      tagArrayWire_18_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_1 <= 22'h0;
    end else if (_T_1460) begin
      tagArrayWire_17_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_1 <= 22'h0;
    end else if (_T_1399) begin
      tagArrayWire_16_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_1 <= 22'h0;
    end else if (_T_1338) begin
      tagArrayWire_15_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_1 <= 22'h0;
    end else if (_T_1277) begin
      tagArrayWire_14_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_1 <= 22'h0;
    end else if (_T_1216) begin
      tagArrayWire_13_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_1 <= 22'h0;
    end else if (_T_1155) begin
      tagArrayWire_12_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_1 <= 22'h0;
    end else if (_T_1094) begin
      tagArrayWire_11_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_1 <= 22'h0;
    end else if (_T_1033) begin
      tagArrayWire_10_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_1 <= 22'h0;
    end else if (_T_972) begin
      tagArrayWire_9_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_1 <= 22'h0;
    end else if (_T_911) begin
      tagArrayWire_8_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_1 <= 22'h0;
    end else if (_T_850) begin
      tagArrayWire_7_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_1 <= 22'h0;
    end else if (_T_789) begin
      tagArrayWire_6_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_1 <= 22'h0;
    end else if (_T_728) begin
      tagArrayWire_5_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_1 <= 22'h0;
    end else if (_T_667) begin
      tagArrayWire_4_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_1 <= 22'h0;
    end else if (_T_606) begin
      tagArrayWire_3_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_1 <= 22'h0;
    end else if (_T_545) begin
      tagArrayWire_2_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_1 <= 22'h0;
    end else if (_T_484) begin
      tagArrayWire_1_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_1 <= 22'h0;
    end else if (_T_423) begin
      tagArrayWire_0_1 <= tag;
    end
    if (_T_412) begin
      vArrayWire_63_2 <= 1'h0;
    end else begin
      vArrayWire_63_2 <= _GEN_573;
    end
    if (_T_412) begin
      vArrayWire_62_2 <= 1'h0;
    end else begin
      vArrayWire_62_2 <= _GEN_564;
    end
    if (_T_412) begin
      vArrayWire_61_2 <= 1'h0;
    end else begin
      vArrayWire_61_2 <= _GEN_555;
    end
    if (_T_412) begin
      vArrayWire_60_2 <= 1'h0;
    end else begin
      vArrayWire_60_2 <= _GEN_546;
    end
    if (_T_412) begin
      vArrayWire_59_2 <= 1'h0;
    end else begin
      vArrayWire_59_2 <= _GEN_537;
    end
    if (_T_412) begin
      vArrayWire_58_2 <= 1'h0;
    end else begin
      vArrayWire_58_2 <= _GEN_528;
    end
    if (_T_412) begin
      vArrayWire_57_2 <= 1'h0;
    end else begin
      vArrayWire_57_2 <= _GEN_519;
    end
    if (_T_412) begin
      vArrayWire_56_2 <= 1'h0;
    end else begin
      vArrayWire_56_2 <= _GEN_510;
    end
    if (_T_412) begin
      vArrayWire_55_2 <= 1'h0;
    end else begin
      vArrayWire_55_2 <= _GEN_501;
    end
    if (_T_412) begin
      vArrayWire_54_2 <= 1'h0;
    end else begin
      vArrayWire_54_2 <= _GEN_492;
    end
    if (_T_412) begin
      vArrayWire_53_2 <= 1'h0;
    end else begin
      vArrayWire_53_2 <= _GEN_483;
    end
    if (_T_412) begin
      vArrayWire_52_2 <= 1'h0;
    end else begin
      vArrayWire_52_2 <= _GEN_474;
    end
    if (_T_412) begin
      vArrayWire_51_2 <= 1'h0;
    end else begin
      vArrayWire_51_2 <= _GEN_465;
    end
    if (_T_412) begin
      vArrayWire_50_2 <= 1'h0;
    end else begin
      vArrayWire_50_2 <= _GEN_456;
    end
    if (_T_412) begin
      vArrayWire_49_2 <= 1'h0;
    end else begin
      vArrayWire_49_2 <= _GEN_447;
    end
    if (_T_412) begin
      vArrayWire_48_2 <= 1'h0;
    end else begin
      vArrayWire_48_2 <= _GEN_438;
    end
    if (_T_412) begin
      vArrayWire_47_2 <= 1'h0;
    end else begin
      vArrayWire_47_2 <= _GEN_429;
    end
    if (_T_412) begin
      vArrayWire_46_2 <= 1'h0;
    end else begin
      vArrayWire_46_2 <= _GEN_420;
    end
    if (_T_412) begin
      vArrayWire_45_2 <= 1'h0;
    end else begin
      vArrayWire_45_2 <= _GEN_411;
    end
    if (_T_412) begin
      vArrayWire_44_2 <= 1'h0;
    end else begin
      vArrayWire_44_2 <= _GEN_402;
    end
    if (_T_412) begin
      vArrayWire_43_2 <= 1'h0;
    end else begin
      vArrayWire_43_2 <= _GEN_393;
    end
    if (_T_412) begin
      vArrayWire_42_2 <= 1'h0;
    end else begin
      vArrayWire_42_2 <= _GEN_384;
    end
    if (_T_412) begin
      vArrayWire_41_2 <= 1'h0;
    end else begin
      vArrayWire_41_2 <= _GEN_375;
    end
    if (_T_412) begin
      vArrayWire_40_2 <= 1'h0;
    end else begin
      vArrayWire_40_2 <= _GEN_366;
    end
    if (_T_412) begin
      vArrayWire_39_2 <= 1'h0;
    end else begin
      vArrayWire_39_2 <= _GEN_357;
    end
    if (_T_412) begin
      vArrayWire_38_2 <= 1'h0;
    end else begin
      vArrayWire_38_2 <= _GEN_348;
    end
    if (_T_412) begin
      vArrayWire_37_2 <= 1'h0;
    end else begin
      vArrayWire_37_2 <= _GEN_339;
    end
    if (_T_412) begin
      vArrayWire_36_2 <= 1'h0;
    end else begin
      vArrayWire_36_2 <= _GEN_330;
    end
    if (_T_412) begin
      vArrayWire_35_2 <= 1'h0;
    end else begin
      vArrayWire_35_2 <= _GEN_321;
    end
    if (_T_412) begin
      vArrayWire_34_2 <= 1'h0;
    end else begin
      vArrayWire_34_2 <= _GEN_312;
    end
    if (_T_412) begin
      vArrayWire_33_2 <= 1'h0;
    end else begin
      vArrayWire_33_2 <= _GEN_303;
    end
    if (_T_412) begin
      vArrayWire_32_2 <= 1'h0;
    end else begin
      vArrayWire_32_2 <= _GEN_294;
    end
    if (_T_412) begin
      vArrayWire_31_2 <= 1'h0;
    end else begin
      vArrayWire_31_2 <= _GEN_285;
    end
    if (_T_412) begin
      vArrayWire_30_2 <= 1'h0;
    end else begin
      vArrayWire_30_2 <= _GEN_276;
    end
    if (_T_412) begin
      vArrayWire_29_2 <= 1'h0;
    end else begin
      vArrayWire_29_2 <= _GEN_267;
    end
    if (_T_412) begin
      vArrayWire_28_2 <= 1'h0;
    end else begin
      vArrayWire_28_2 <= _GEN_258;
    end
    if (_T_412) begin
      vArrayWire_27_2 <= 1'h0;
    end else begin
      vArrayWire_27_2 <= _GEN_249;
    end
    if (_T_412) begin
      vArrayWire_26_2 <= 1'h0;
    end else begin
      vArrayWire_26_2 <= _GEN_240;
    end
    if (_T_412) begin
      vArrayWire_25_2 <= 1'h0;
    end else begin
      vArrayWire_25_2 <= _GEN_231;
    end
    if (_T_412) begin
      vArrayWire_24_2 <= 1'h0;
    end else begin
      vArrayWire_24_2 <= _GEN_222;
    end
    if (_T_412) begin
      vArrayWire_23_2 <= 1'h0;
    end else begin
      vArrayWire_23_2 <= _GEN_213;
    end
    if (_T_412) begin
      vArrayWire_22_2 <= 1'h0;
    end else begin
      vArrayWire_22_2 <= _GEN_204;
    end
    if (_T_412) begin
      vArrayWire_21_2 <= 1'h0;
    end else begin
      vArrayWire_21_2 <= _GEN_195;
    end
    if (_T_412) begin
      vArrayWire_20_2 <= 1'h0;
    end else begin
      vArrayWire_20_2 <= _GEN_186;
    end
    if (_T_412) begin
      vArrayWire_19_2 <= 1'h0;
    end else begin
      vArrayWire_19_2 <= _GEN_177;
    end
    if (_T_412) begin
      vArrayWire_18_2 <= 1'h0;
    end else begin
      vArrayWire_18_2 <= _GEN_168;
    end
    if (_T_412) begin
      vArrayWire_17_2 <= 1'h0;
    end else begin
      vArrayWire_17_2 <= _GEN_159;
    end
    if (_T_412) begin
      vArrayWire_16_2 <= 1'h0;
    end else begin
      vArrayWire_16_2 <= _GEN_150;
    end
    if (_T_412) begin
      vArrayWire_15_2 <= 1'h0;
    end else begin
      vArrayWire_15_2 <= _GEN_141;
    end
    if (_T_412) begin
      vArrayWire_14_2 <= 1'h0;
    end else begin
      vArrayWire_14_2 <= _GEN_132;
    end
    if (_T_412) begin
      vArrayWire_13_2 <= 1'h0;
    end else begin
      vArrayWire_13_2 <= _GEN_123;
    end
    if (_T_412) begin
      vArrayWire_12_2 <= 1'h0;
    end else begin
      vArrayWire_12_2 <= _GEN_114;
    end
    if (_T_412) begin
      vArrayWire_11_2 <= 1'h0;
    end else begin
      vArrayWire_11_2 <= _GEN_105;
    end
    if (_T_412) begin
      vArrayWire_10_2 <= 1'h0;
    end else begin
      vArrayWire_10_2 <= _GEN_96;
    end
    if (_T_412) begin
      vArrayWire_9_2 <= 1'h0;
    end else begin
      vArrayWire_9_2 <= _GEN_87;
    end
    if (_T_412) begin
      vArrayWire_8_2 <= 1'h0;
    end else begin
      vArrayWire_8_2 <= _GEN_78;
    end
    if (_T_412) begin
      vArrayWire_7_2 <= 1'h0;
    end else begin
      vArrayWire_7_2 <= _GEN_69;
    end
    if (_T_412) begin
      vArrayWire_6_2 <= 1'h0;
    end else begin
      vArrayWire_6_2 <= _GEN_60;
    end
    if (_T_412) begin
      vArrayWire_5_2 <= 1'h0;
    end else begin
      vArrayWire_5_2 <= _GEN_51;
    end
    if (_T_412) begin
      vArrayWire_4_2 <= 1'h0;
    end else begin
      vArrayWire_4_2 <= _GEN_42;
    end
    if (_T_412) begin
      vArrayWire_3_2 <= 1'h0;
    end else begin
      vArrayWire_3_2 <= _GEN_33;
    end
    if (_T_412) begin
      vArrayWire_2_2 <= 1'h0;
    end else begin
      vArrayWire_2_2 <= _GEN_24;
    end
    if (_T_412) begin
      vArrayWire_1_2 <= 1'h0;
    end else begin
      vArrayWire_1_2 <= _GEN_15;
    end
    if (_T_412) begin
      vArrayWire_0_2 <= 1'h0;
    end else begin
      vArrayWire_0_2 <= _GEN_6;
    end
    if (reset) begin
      tagArrayWire_63_2 <= 22'h0;
    end else if (_T_4280) begin
      tagArrayWire_63_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_2 <= 22'h0;
    end else if (_T_4219) begin
      tagArrayWire_62_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_2 <= 22'h0;
    end else if (_T_4158) begin
      tagArrayWire_61_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_2 <= 22'h0;
    end else if (_T_4097) begin
      tagArrayWire_60_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_2 <= 22'h0;
    end else if (_T_4036) begin
      tagArrayWire_59_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_2 <= 22'h0;
    end else if (_T_3975) begin
      tagArrayWire_58_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_2 <= 22'h0;
    end else if (_T_3914) begin
      tagArrayWire_57_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_2 <= 22'h0;
    end else if (_T_3853) begin
      tagArrayWire_56_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_2 <= 22'h0;
    end else if (_T_3792) begin
      tagArrayWire_55_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_2 <= 22'h0;
    end else if (_T_3731) begin
      tagArrayWire_54_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_2 <= 22'h0;
    end else if (_T_3670) begin
      tagArrayWire_53_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_2 <= 22'h0;
    end else if (_T_3609) begin
      tagArrayWire_52_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_2 <= 22'h0;
    end else if (_T_3548) begin
      tagArrayWire_51_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_2 <= 22'h0;
    end else if (_T_3487) begin
      tagArrayWire_50_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_2 <= 22'h0;
    end else if (_T_3426) begin
      tagArrayWire_49_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_2 <= 22'h0;
    end else if (_T_3365) begin
      tagArrayWire_48_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_2 <= 22'h0;
    end else if (_T_3304) begin
      tagArrayWire_47_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_2 <= 22'h0;
    end else if (_T_3243) begin
      tagArrayWire_46_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_2 <= 22'h0;
    end else if (_T_3182) begin
      tagArrayWire_45_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_2 <= 22'h0;
    end else if (_T_3121) begin
      tagArrayWire_44_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_2 <= 22'h0;
    end else if (_T_3060) begin
      tagArrayWire_43_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_2 <= 22'h0;
    end else if (_T_2999) begin
      tagArrayWire_42_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_2 <= 22'h0;
    end else if (_T_2938) begin
      tagArrayWire_41_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_2 <= 22'h0;
    end else if (_T_2877) begin
      tagArrayWire_40_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_2 <= 22'h0;
    end else if (_T_2816) begin
      tagArrayWire_39_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_2 <= 22'h0;
    end else if (_T_2755) begin
      tagArrayWire_38_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_2 <= 22'h0;
    end else if (_T_2694) begin
      tagArrayWire_37_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_2 <= 22'h0;
    end else if (_T_2633) begin
      tagArrayWire_36_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_2 <= 22'h0;
    end else if (_T_2572) begin
      tagArrayWire_35_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_2 <= 22'h0;
    end else if (_T_2511) begin
      tagArrayWire_34_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_2 <= 22'h0;
    end else if (_T_2450) begin
      tagArrayWire_33_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_2 <= 22'h0;
    end else if (_T_2389) begin
      tagArrayWire_32_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_2 <= 22'h0;
    end else if (_T_2328) begin
      tagArrayWire_31_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_2 <= 22'h0;
    end else if (_T_2267) begin
      tagArrayWire_30_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_2 <= 22'h0;
    end else if (_T_2206) begin
      tagArrayWire_29_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_2 <= 22'h0;
    end else if (_T_2145) begin
      tagArrayWire_28_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_2 <= 22'h0;
    end else if (_T_2084) begin
      tagArrayWire_27_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_2 <= 22'h0;
    end else if (_T_2023) begin
      tagArrayWire_26_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_2 <= 22'h0;
    end else if (_T_1962) begin
      tagArrayWire_25_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_2 <= 22'h0;
    end else if (_T_1901) begin
      tagArrayWire_24_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_2 <= 22'h0;
    end else if (_T_1840) begin
      tagArrayWire_23_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_2 <= 22'h0;
    end else if (_T_1779) begin
      tagArrayWire_22_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_2 <= 22'h0;
    end else if (_T_1718) begin
      tagArrayWire_21_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_2 <= 22'h0;
    end else if (_T_1657) begin
      tagArrayWire_20_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_2 <= 22'h0;
    end else if (_T_1596) begin
      tagArrayWire_19_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_2 <= 22'h0;
    end else if (_T_1535) begin
      tagArrayWire_18_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_2 <= 22'h0;
    end else if (_T_1474) begin
      tagArrayWire_17_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_2 <= 22'h0;
    end else if (_T_1413) begin
      tagArrayWire_16_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_2 <= 22'h0;
    end else if (_T_1352) begin
      tagArrayWire_15_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_2 <= 22'h0;
    end else if (_T_1291) begin
      tagArrayWire_14_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_2 <= 22'h0;
    end else if (_T_1230) begin
      tagArrayWire_13_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_2 <= 22'h0;
    end else if (_T_1169) begin
      tagArrayWire_12_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_2 <= 22'h0;
    end else if (_T_1108) begin
      tagArrayWire_11_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_2 <= 22'h0;
    end else if (_T_1047) begin
      tagArrayWire_10_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_2 <= 22'h0;
    end else if (_T_986) begin
      tagArrayWire_9_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_2 <= 22'h0;
    end else if (_T_925) begin
      tagArrayWire_8_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_2 <= 22'h0;
    end else if (_T_864) begin
      tagArrayWire_7_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_2 <= 22'h0;
    end else if (_T_803) begin
      tagArrayWire_6_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_2 <= 22'h0;
    end else if (_T_742) begin
      tagArrayWire_5_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_2 <= 22'h0;
    end else if (_T_681) begin
      tagArrayWire_4_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_2 <= 22'h0;
    end else if (_T_620) begin
      tagArrayWire_3_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_2 <= 22'h0;
    end else if (_T_559) begin
      tagArrayWire_2_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_2 <= 22'h0;
    end else if (_T_498) begin
      tagArrayWire_1_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_2 <= 22'h0;
    end else if (_T_437) begin
      tagArrayWire_0_2 <= tag;
    end
    if (_T_412) begin
      vArrayWire_63_3 <= 1'h0;
    end else begin
      vArrayWire_63_3 <= _GEN_575;
    end
    if (_T_412) begin
      vArrayWire_62_3 <= 1'h0;
    end else begin
      vArrayWire_62_3 <= _GEN_566;
    end
    if (_T_412) begin
      vArrayWire_61_3 <= 1'h0;
    end else begin
      vArrayWire_61_3 <= _GEN_557;
    end
    if (_T_412) begin
      vArrayWire_60_3 <= 1'h0;
    end else begin
      vArrayWire_60_3 <= _GEN_548;
    end
    if (_T_412) begin
      vArrayWire_59_3 <= 1'h0;
    end else begin
      vArrayWire_59_3 <= _GEN_539;
    end
    if (_T_412) begin
      vArrayWire_58_3 <= 1'h0;
    end else begin
      vArrayWire_58_3 <= _GEN_530;
    end
    if (_T_412) begin
      vArrayWire_57_3 <= 1'h0;
    end else begin
      vArrayWire_57_3 <= _GEN_521;
    end
    if (_T_412) begin
      vArrayWire_56_3 <= 1'h0;
    end else begin
      vArrayWire_56_3 <= _GEN_512;
    end
    if (_T_412) begin
      vArrayWire_55_3 <= 1'h0;
    end else begin
      vArrayWire_55_3 <= _GEN_503;
    end
    if (_T_412) begin
      vArrayWire_54_3 <= 1'h0;
    end else begin
      vArrayWire_54_3 <= _GEN_494;
    end
    if (_T_412) begin
      vArrayWire_53_3 <= 1'h0;
    end else begin
      vArrayWire_53_3 <= _GEN_485;
    end
    if (_T_412) begin
      vArrayWire_52_3 <= 1'h0;
    end else begin
      vArrayWire_52_3 <= _GEN_476;
    end
    if (_T_412) begin
      vArrayWire_51_3 <= 1'h0;
    end else begin
      vArrayWire_51_3 <= _GEN_467;
    end
    if (_T_412) begin
      vArrayWire_50_3 <= 1'h0;
    end else begin
      vArrayWire_50_3 <= _GEN_458;
    end
    if (_T_412) begin
      vArrayWire_49_3 <= 1'h0;
    end else begin
      vArrayWire_49_3 <= _GEN_449;
    end
    if (_T_412) begin
      vArrayWire_48_3 <= 1'h0;
    end else begin
      vArrayWire_48_3 <= _GEN_440;
    end
    if (_T_412) begin
      vArrayWire_47_3 <= 1'h0;
    end else begin
      vArrayWire_47_3 <= _GEN_431;
    end
    if (_T_412) begin
      vArrayWire_46_3 <= 1'h0;
    end else begin
      vArrayWire_46_3 <= _GEN_422;
    end
    if (_T_412) begin
      vArrayWire_45_3 <= 1'h0;
    end else begin
      vArrayWire_45_3 <= _GEN_413;
    end
    if (_T_412) begin
      vArrayWire_44_3 <= 1'h0;
    end else begin
      vArrayWire_44_3 <= _GEN_404;
    end
    if (_T_412) begin
      vArrayWire_43_3 <= 1'h0;
    end else begin
      vArrayWire_43_3 <= _GEN_395;
    end
    if (_T_412) begin
      vArrayWire_42_3 <= 1'h0;
    end else begin
      vArrayWire_42_3 <= _GEN_386;
    end
    if (_T_412) begin
      vArrayWire_41_3 <= 1'h0;
    end else begin
      vArrayWire_41_3 <= _GEN_377;
    end
    if (_T_412) begin
      vArrayWire_40_3 <= 1'h0;
    end else begin
      vArrayWire_40_3 <= _GEN_368;
    end
    if (_T_412) begin
      vArrayWire_39_3 <= 1'h0;
    end else begin
      vArrayWire_39_3 <= _GEN_359;
    end
    if (_T_412) begin
      vArrayWire_38_3 <= 1'h0;
    end else begin
      vArrayWire_38_3 <= _GEN_350;
    end
    if (_T_412) begin
      vArrayWire_37_3 <= 1'h0;
    end else begin
      vArrayWire_37_3 <= _GEN_341;
    end
    if (_T_412) begin
      vArrayWire_36_3 <= 1'h0;
    end else begin
      vArrayWire_36_3 <= _GEN_332;
    end
    if (_T_412) begin
      vArrayWire_35_3 <= 1'h0;
    end else begin
      vArrayWire_35_3 <= _GEN_323;
    end
    if (_T_412) begin
      vArrayWire_34_3 <= 1'h0;
    end else begin
      vArrayWire_34_3 <= _GEN_314;
    end
    if (_T_412) begin
      vArrayWire_33_3 <= 1'h0;
    end else begin
      vArrayWire_33_3 <= _GEN_305;
    end
    if (_T_412) begin
      vArrayWire_32_3 <= 1'h0;
    end else begin
      vArrayWire_32_3 <= _GEN_296;
    end
    if (_T_412) begin
      vArrayWire_31_3 <= 1'h0;
    end else begin
      vArrayWire_31_3 <= _GEN_287;
    end
    if (_T_412) begin
      vArrayWire_30_3 <= 1'h0;
    end else begin
      vArrayWire_30_3 <= _GEN_278;
    end
    if (_T_412) begin
      vArrayWire_29_3 <= 1'h0;
    end else begin
      vArrayWire_29_3 <= _GEN_269;
    end
    if (_T_412) begin
      vArrayWire_28_3 <= 1'h0;
    end else begin
      vArrayWire_28_3 <= _GEN_260;
    end
    if (_T_412) begin
      vArrayWire_27_3 <= 1'h0;
    end else begin
      vArrayWire_27_3 <= _GEN_251;
    end
    if (_T_412) begin
      vArrayWire_26_3 <= 1'h0;
    end else begin
      vArrayWire_26_3 <= _GEN_242;
    end
    if (_T_412) begin
      vArrayWire_25_3 <= 1'h0;
    end else begin
      vArrayWire_25_3 <= _GEN_233;
    end
    if (_T_412) begin
      vArrayWire_24_3 <= 1'h0;
    end else begin
      vArrayWire_24_3 <= _GEN_224;
    end
    if (_T_412) begin
      vArrayWire_23_3 <= 1'h0;
    end else begin
      vArrayWire_23_3 <= _GEN_215;
    end
    if (_T_412) begin
      vArrayWire_22_3 <= 1'h0;
    end else begin
      vArrayWire_22_3 <= _GEN_206;
    end
    if (_T_412) begin
      vArrayWire_21_3 <= 1'h0;
    end else begin
      vArrayWire_21_3 <= _GEN_197;
    end
    if (_T_412) begin
      vArrayWire_20_3 <= 1'h0;
    end else begin
      vArrayWire_20_3 <= _GEN_188;
    end
    if (_T_412) begin
      vArrayWire_19_3 <= 1'h0;
    end else begin
      vArrayWire_19_3 <= _GEN_179;
    end
    if (_T_412) begin
      vArrayWire_18_3 <= 1'h0;
    end else begin
      vArrayWire_18_3 <= _GEN_170;
    end
    if (_T_412) begin
      vArrayWire_17_3 <= 1'h0;
    end else begin
      vArrayWire_17_3 <= _GEN_161;
    end
    if (_T_412) begin
      vArrayWire_16_3 <= 1'h0;
    end else begin
      vArrayWire_16_3 <= _GEN_152;
    end
    if (_T_412) begin
      vArrayWire_15_3 <= 1'h0;
    end else begin
      vArrayWire_15_3 <= _GEN_143;
    end
    if (_T_412) begin
      vArrayWire_14_3 <= 1'h0;
    end else begin
      vArrayWire_14_3 <= _GEN_134;
    end
    if (_T_412) begin
      vArrayWire_13_3 <= 1'h0;
    end else begin
      vArrayWire_13_3 <= _GEN_125;
    end
    if (_T_412) begin
      vArrayWire_12_3 <= 1'h0;
    end else begin
      vArrayWire_12_3 <= _GEN_116;
    end
    if (_T_412) begin
      vArrayWire_11_3 <= 1'h0;
    end else begin
      vArrayWire_11_3 <= _GEN_107;
    end
    if (_T_412) begin
      vArrayWire_10_3 <= 1'h0;
    end else begin
      vArrayWire_10_3 <= _GEN_98;
    end
    if (_T_412) begin
      vArrayWire_9_3 <= 1'h0;
    end else begin
      vArrayWire_9_3 <= _GEN_89;
    end
    if (_T_412) begin
      vArrayWire_8_3 <= 1'h0;
    end else begin
      vArrayWire_8_3 <= _GEN_80;
    end
    if (_T_412) begin
      vArrayWire_7_3 <= 1'h0;
    end else begin
      vArrayWire_7_3 <= _GEN_71;
    end
    if (_T_412) begin
      vArrayWire_6_3 <= 1'h0;
    end else begin
      vArrayWire_6_3 <= _GEN_62;
    end
    if (_T_412) begin
      vArrayWire_5_3 <= 1'h0;
    end else begin
      vArrayWire_5_3 <= _GEN_53;
    end
    if (_T_412) begin
      vArrayWire_4_3 <= 1'h0;
    end else begin
      vArrayWire_4_3 <= _GEN_44;
    end
    if (_T_412) begin
      vArrayWire_3_3 <= 1'h0;
    end else begin
      vArrayWire_3_3 <= _GEN_35;
    end
    if (_T_412) begin
      vArrayWire_2_3 <= 1'h0;
    end else begin
      vArrayWire_2_3 <= _GEN_26;
    end
    if (_T_412) begin
      vArrayWire_1_3 <= 1'h0;
    end else begin
      vArrayWire_1_3 <= _GEN_17;
    end
    if (_T_412) begin
      vArrayWire_0_3 <= 1'h0;
    end else begin
      vArrayWire_0_3 <= _GEN_8;
    end
    if (reset) begin
      tagArrayWire_63_3 <= 22'h0;
    end else if (_T_4294) begin
      tagArrayWire_63_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_3 <= 22'h0;
    end else if (_T_4233) begin
      tagArrayWire_62_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_3 <= 22'h0;
    end else if (_T_4172) begin
      tagArrayWire_61_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_3 <= 22'h0;
    end else if (_T_4111) begin
      tagArrayWire_60_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_3 <= 22'h0;
    end else if (_T_4050) begin
      tagArrayWire_59_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_3 <= 22'h0;
    end else if (_T_3989) begin
      tagArrayWire_58_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_3 <= 22'h0;
    end else if (_T_3928) begin
      tagArrayWire_57_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_3 <= 22'h0;
    end else if (_T_3867) begin
      tagArrayWire_56_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_3 <= 22'h0;
    end else if (_T_3806) begin
      tagArrayWire_55_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_3 <= 22'h0;
    end else if (_T_3745) begin
      tagArrayWire_54_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_3 <= 22'h0;
    end else if (_T_3684) begin
      tagArrayWire_53_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_3 <= 22'h0;
    end else if (_T_3623) begin
      tagArrayWire_52_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_3 <= 22'h0;
    end else if (_T_3562) begin
      tagArrayWire_51_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_3 <= 22'h0;
    end else if (_T_3501) begin
      tagArrayWire_50_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_3 <= 22'h0;
    end else if (_T_3440) begin
      tagArrayWire_49_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_3 <= 22'h0;
    end else if (_T_3379) begin
      tagArrayWire_48_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_3 <= 22'h0;
    end else if (_T_3318) begin
      tagArrayWire_47_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_3 <= 22'h0;
    end else if (_T_3257) begin
      tagArrayWire_46_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_3 <= 22'h0;
    end else if (_T_3196) begin
      tagArrayWire_45_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_3 <= 22'h0;
    end else if (_T_3135) begin
      tagArrayWire_44_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_3 <= 22'h0;
    end else if (_T_3074) begin
      tagArrayWire_43_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_3 <= 22'h0;
    end else if (_T_3013) begin
      tagArrayWire_42_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_3 <= 22'h0;
    end else if (_T_2952) begin
      tagArrayWire_41_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_3 <= 22'h0;
    end else if (_T_2891) begin
      tagArrayWire_40_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_3 <= 22'h0;
    end else if (_T_2830) begin
      tagArrayWire_39_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_3 <= 22'h0;
    end else if (_T_2769) begin
      tagArrayWire_38_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_3 <= 22'h0;
    end else if (_T_2708) begin
      tagArrayWire_37_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_3 <= 22'h0;
    end else if (_T_2647) begin
      tagArrayWire_36_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_3 <= 22'h0;
    end else if (_T_2586) begin
      tagArrayWire_35_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_3 <= 22'h0;
    end else if (_T_2525) begin
      tagArrayWire_34_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_3 <= 22'h0;
    end else if (_T_2464) begin
      tagArrayWire_33_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_3 <= 22'h0;
    end else if (_T_2403) begin
      tagArrayWire_32_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_3 <= 22'h0;
    end else if (_T_2342) begin
      tagArrayWire_31_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_3 <= 22'h0;
    end else if (_T_2281) begin
      tagArrayWire_30_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_3 <= 22'h0;
    end else if (_T_2220) begin
      tagArrayWire_29_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_3 <= 22'h0;
    end else if (_T_2159) begin
      tagArrayWire_28_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_3 <= 22'h0;
    end else if (_T_2098) begin
      tagArrayWire_27_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_3 <= 22'h0;
    end else if (_T_2037) begin
      tagArrayWire_26_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_3 <= 22'h0;
    end else if (_T_1976) begin
      tagArrayWire_25_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_3 <= 22'h0;
    end else if (_T_1915) begin
      tagArrayWire_24_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_3 <= 22'h0;
    end else if (_T_1854) begin
      tagArrayWire_23_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_3 <= 22'h0;
    end else if (_T_1793) begin
      tagArrayWire_22_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_3 <= 22'h0;
    end else if (_T_1732) begin
      tagArrayWire_21_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_3 <= 22'h0;
    end else if (_T_1671) begin
      tagArrayWire_20_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_3 <= 22'h0;
    end else if (_T_1610) begin
      tagArrayWire_19_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_3 <= 22'h0;
    end else if (_T_1549) begin
      tagArrayWire_18_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_3 <= 22'h0;
    end else if (_T_1488) begin
      tagArrayWire_17_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_3 <= 22'h0;
    end else if (_T_1427) begin
      tagArrayWire_16_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_3 <= 22'h0;
    end else if (_T_1366) begin
      tagArrayWire_15_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_3 <= 22'h0;
    end else if (_T_1305) begin
      tagArrayWire_14_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_3 <= 22'h0;
    end else if (_T_1244) begin
      tagArrayWire_13_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_3 <= 22'h0;
    end else if (_T_1183) begin
      tagArrayWire_12_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_3 <= 22'h0;
    end else if (_T_1122) begin
      tagArrayWire_11_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_3 <= 22'h0;
    end else if (_T_1061) begin
      tagArrayWire_10_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_3 <= 22'h0;
    end else if (_T_1000) begin
      tagArrayWire_9_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_3 <= 22'h0;
    end else if (_T_939) begin
      tagArrayWire_8_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_3 <= 22'h0;
    end else if (_T_878) begin
      tagArrayWire_7_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_3 <= 22'h0;
    end else if (_T_817) begin
      tagArrayWire_6_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_3 <= 22'h0;
    end else if (_T_756) begin
      tagArrayWire_5_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_3 <= 22'h0;
    end else if (_T_695) begin
      tagArrayWire_4_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_3 <= 22'h0;
    end else if (_T_634) begin
      tagArrayWire_3_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_3 <= 22'h0;
    end else if (_T_573) begin
      tagArrayWire_2_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_3 <= 22'h0;
    end else if (_T_512) begin
      tagArrayWire_1_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_3 <= 22'h0;
    end else if (_T_451) begin
      tagArrayWire_0_3 <= tag;
    end
    if (reset) begin
      selArrayWire_1 <= 2'h0;
    end else if (_T_464) begin
      selArrayWire_1 <= _T_462;
    end
    if (reset) begin
      selArrayWire_0 <= 2'h0;
    end else if (_T_403) begin
      selArrayWire_0 <= _T_401;
    end
    if (reset) begin
      selArrayWire_2 <= 2'h0;
    end else if (_T_525) begin
      selArrayWire_2 <= _T_523;
    end
    if (reset) begin
      selArrayWire_3 <= 2'h0;
    end else if (_T_586) begin
      selArrayWire_3 <= _T_584;
    end
    if (reset) begin
      selArrayWire_4 <= 2'h0;
    end else if (_T_647) begin
      selArrayWire_4 <= _T_645;
    end
    if (reset) begin
      selArrayWire_5 <= 2'h0;
    end else if (_T_708) begin
      selArrayWire_5 <= _T_706;
    end
    if (reset) begin
      selArrayWire_6 <= 2'h0;
    end else if (_T_769) begin
      selArrayWire_6 <= _T_767;
    end
    if (reset) begin
      selArrayWire_7 <= 2'h0;
    end else if (_T_830) begin
      selArrayWire_7 <= _T_828;
    end
    if (reset) begin
      selArrayWire_8 <= 2'h0;
    end else if (_T_891) begin
      selArrayWire_8 <= _T_889;
    end
    if (reset) begin
      selArrayWire_9 <= 2'h0;
    end else if (_T_952) begin
      selArrayWire_9 <= _T_950;
    end
    if (reset) begin
      selArrayWire_10 <= 2'h0;
    end else if (_T_1013) begin
      selArrayWire_10 <= _T_1011;
    end
    if (reset) begin
      selArrayWire_11 <= 2'h0;
    end else if (_T_1074) begin
      selArrayWire_11 <= _T_1072;
    end
    if (reset) begin
      selArrayWire_12 <= 2'h0;
    end else if (_T_1135) begin
      selArrayWire_12 <= _T_1133;
    end
    if (reset) begin
      selArrayWire_13 <= 2'h0;
    end else if (_T_1196) begin
      selArrayWire_13 <= _T_1194;
    end
    if (reset) begin
      selArrayWire_14 <= 2'h0;
    end else if (_T_1257) begin
      selArrayWire_14 <= _T_1255;
    end
    if (reset) begin
      selArrayWire_15 <= 2'h0;
    end else if (_T_1318) begin
      selArrayWire_15 <= _T_1316;
    end
    if (reset) begin
      selArrayWire_16 <= 2'h0;
    end else if (_T_1379) begin
      selArrayWire_16 <= _T_1377;
    end
    if (reset) begin
      selArrayWire_17 <= 2'h0;
    end else if (_T_1440) begin
      selArrayWire_17 <= _T_1438;
    end
    if (reset) begin
      selArrayWire_18 <= 2'h0;
    end else if (_T_1501) begin
      selArrayWire_18 <= _T_1499;
    end
    if (reset) begin
      selArrayWire_19 <= 2'h0;
    end else if (_T_1562) begin
      selArrayWire_19 <= _T_1560;
    end
    if (reset) begin
      selArrayWire_20 <= 2'h0;
    end else if (_T_1623) begin
      selArrayWire_20 <= _T_1621;
    end
    if (reset) begin
      selArrayWire_21 <= 2'h0;
    end else if (_T_1684) begin
      selArrayWire_21 <= _T_1682;
    end
    if (reset) begin
      selArrayWire_22 <= 2'h0;
    end else if (_T_1745) begin
      selArrayWire_22 <= _T_1743;
    end
    if (reset) begin
      selArrayWire_23 <= 2'h0;
    end else if (_T_1806) begin
      selArrayWire_23 <= _T_1804;
    end
    if (reset) begin
      selArrayWire_24 <= 2'h0;
    end else if (_T_1867) begin
      selArrayWire_24 <= _T_1865;
    end
    if (reset) begin
      selArrayWire_25 <= 2'h0;
    end else if (_T_1928) begin
      selArrayWire_25 <= _T_1926;
    end
    if (reset) begin
      selArrayWire_26 <= 2'h0;
    end else if (_T_1989) begin
      selArrayWire_26 <= _T_1987;
    end
    if (reset) begin
      selArrayWire_27 <= 2'h0;
    end else if (_T_2050) begin
      selArrayWire_27 <= _T_2048;
    end
    if (reset) begin
      selArrayWire_28 <= 2'h0;
    end else if (_T_2111) begin
      selArrayWire_28 <= _T_2109;
    end
    if (reset) begin
      selArrayWire_29 <= 2'h0;
    end else if (_T_2172) begin
      selArrayWire_29 <= _T_2170;
    end
    if (reset) begin
      selArrayWire_30 <= 2'h0;
    end else if (_T_2233) begin
      selArrayWire_30 <= _T_2231;
    end
    if (reset) begin
      selArrayWire_31 <= 2'h0;
    end else if (_T_2294) begin
      selArrayWire_31 <= _T_2292;
    end
    if (reset) begin
      selArrayWire_32 <= 2'h0;
    end else if (_T_2355) begin
      selArrayWire_32 <= _T_2353;
    end
    if (reset) begin
      selArrayWire_33 <= 2'h0;
    end else if (_T_2416) begin
      selArrayWire_33 <= _T_2414;
    end
    if (reset) begin
      selArrayWire_34 <= 2'h0;
    end else if (_T_2477) begin
      selArrayWire_34 <= _T_2475;
    end
    if (reset) begin
      selArrayWire_35 <= 2'h0;
    end else if (_T_2538) begin
      selArrayWire_35 <= _T_2536;
    end
    if (reset) begin
      selArrayWire_36 <= 2'h0;
    end else if (_T_2599) begin
      selArrayWire_36 <= _T_2597;
    end
    if (reset) begin
      selArrayWire_37 <= 2'h0;
    end else if (_T_2660) begin
      selArrayWire_37 <= _T_2658;
    end
    if (reset) begin
      selArrayWire_38 <= 2'h0;
    end else if (_T_2721) begin
      selArrayWire_38 <= _T_2719;
    end
    if (reset) begin
      selArrayWire_39 <= 2'h0;
    end else if (_T_2782) begin
      selArrayWire_39 <= _T_2780;
    end
    if (reset) begin
      selArrayWire_40 <= 2'h0;
    end else if (_T_2843) begin
      selArrayWire_40 <= _T_2841;
    end
    if (reset) begin
      selArrayWire_41 <= 2'h0;
    end else if (_T_2904) begin
      selArrayWire_41 <= _T_2902;
    end
    if (reset) begin
      selArrayWire_42 <= 2'h0;
    end else if (_T_2965) begin
      selArrayWire_42 <= _T_2963;
    end
    if (reset) begin
      selArrayWire_43 <= 2'h0;
    end else if (_T_3026) begin
      selArrayWire_43 <= _T_3024;
    end
    if (reset) begin
      selArrayWire_44 <= 2'h0;
    end else if (_T_3087) begin
      selArrayWire_44 <= _T_3085;
    end
    if (reset) begin
      selArrayWire_45 <= 2'h0;
    end else if (_T_3148) begin
      selArrayWire_45 <= _T_3146;
    end
    if (reset) begin
      selArrayWire_46 <= 2'h0;
    end else if (_T_3209) begin
      selArrayWire_46 <= _T_3207;
    end
    if (reset) begin
      selArrayWire_47 <= 2'h0;
    end else if (_T_3270) begin
      selArrayWire_47 <= _T_3268;
    end
    if (reset) begin
      selArrayWire_48 <= 2'h0;
    end else if (_T_3331) begin
      selArrayWire_48 <= _T_3329;
    end
    if (reset) begin
      selArrayWire_49 <= 2'h0;
    end else if (_T_3392) begin
      selArrayWire_49 <= _T_3390;
    end
    if (reset) begin
      selArrayWire_50 <= 2'h0;
    end else if (_T_3453) begin
      selArrayWire_50 <= _T_3451;
    end
    if (reset) begin
      selArrayWire_51 <= 2'h0;
    end else if (_T_3514) begin
      selArrayWire_51 <= _T_3512;
    end
    if (reset) begin
      selArrayWire_52 <= 2'h0;
    end else if (_T_3575) begin
      selArrayWire_52 <= _T_3573;
    end
    if (reset) begin
      selArrayWire_53 <= 2'h0;
    end else if (_T_3636) begin
      selArrayWire_53 <= _T_3634;
    end
    if (reset) begin
      selArrayWire_54 <= 2'h0;
    end else if (_T_3697) begin
      selArrayWire_54 <= _T_3695;
    end
    if (reset) begin
      selArrayWire_55 <= 2'h0;
    end else if (_T_3758) begin
      selArrayWire_55 <= _T_3756;
    end
    if (reset) begin
      selArrayWire_56 <= 2'h0;
    end else if (_T_3819) begin
      selArrayWire_56 <= _T_3817;
    end
    if (reset) begin
      selArrayWire_57 <= 2'h0;
    end else if (_T_3880) begin
      selArrayWire_57 <= _T_3878;
    end
    if (reset) begin
      selArrayWire_58 <= 2'h0;
    end else if (_T_3941) begin
      selArrayWire_58 <= _T_3939;
    end
    if (reset) begin
      selArrayWire_59 <= 2'h0;
    end else if (_T_4002) begin
      selArrayWire_59 <= _T_4000;
    end
    if (reset) begin
      selArrayWire_60 <= 2'h0;
    end else if (_T_4063) begin
      selArrayWire_60 <= _T_4061;
    end
    if (reset) begin
      selArrayWire_61 <= 2'h0;
    end else if (_T_4124) begin
      selArrayWire_61 <= _T_4122;
    end
    if (reset) begin
      selArrayWire_62 <= 2'h0;
    end else if (_T_4185) begin
      selArrayWire_62 <= _T_4183;
    end
    if (reset) begin
      selArrayWire_63 <= 2'h0;
    end else if (_T_4246) begin
      selArrayWire_63 <= _T_4244;
    end
  end
endmodule
module AXICache(
  input         clock,
  input         reset,
  input         io_axiIO_awready,
  output        io_axiIO_awvalid,
  output [31:0] io_axiIO_awaddr,
  output [2:0]  io_axiIO_awsize,
  input         io_axiIO_wready,
  output        io_axiIO_wvalid,
  output [63:0] io_axiIO_wdata,
  output [7:0]  io_axiIO_wstrb,
  output        io_axiIO_wlast,
  output        io_axiIO_bready,
  input         io_axiIO_bvalid,
  input         io_axiIO_arready,
  output        io_axiIO_arvalid,
  output [31:0] io_axiIO_araddr,
  output [7:0]  io_axiIO_arlen,
  output [2:0]  io_axiIO_arsize,
  output [1:0]  io_axiIO_arburst,
  output        io_axiIO_rready,
  input         io_axiIO_rvalid,
  input  [63:0] io_axiIO_rdata,
  input         io_axiIO_rlast,
  input         io_cache_ar_valid_o,
  input  [31:0] io_cache_ar_addr_o,
  input  [7:0]  io_cache_ar_len_o,
  output        io_cache_r_valid_i,
  output [63:0] io_cache_r_data_i,
  output        io_cache_r_last_i,
  input         io_cache_w_valid_o,
  output        io_cache_w_ready_i,
  input  [63:0] io_cache_w_data_o,
  input  [31:0] io_cache_w_addr_o,
  input  [7:0]  io_cache_w_mask_o,
  input  [1:0]  io_cache_wsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rd_state; // @[AXICache.scala 25:25]
  wire  _T = io_axiIO_rlast & io_axiIO_rvalid; // @[AXICache.scala 30:22]
  wire  _T_3 = 2'h0 == rd_state; // @[Mux.scala 80:60]
  wire  _T_5 = 2'h1 == rd_state; // @[Mux.scala 80:60]
  wire  _T_7 = 2'h2 == rd_state; // @[Mux.scala 80:60]
  wire  isReq = rd_state == 2'h1; // @[AXICache.scala 46:24]
  wire  isData = rd_state == 2'h2; // @[AXICache.scala 47:25]
  wire [1:0] _T_12 = isReq ? 2'h3 : 2'h0; // @[AXICache.scala 62:25]
  wire [1:0] valid_c = {io_axiIO_awready,io_axiIO_wready}; // @[Cat.scala 29:58]
  reg [1:0] w_state; // @[AXICache.scala 75:24]
  wire  _T_15 = 2'h2 == valid_c; // @[Mux.scala 80:60]
  wire  _T_17 = 2'h3 == valid_c; // @[Mux.scala 80:60]
  wire  _T_18 = 2'h1 == w_state; // @[Mux.scala 80:60]
  wire  _T_20 = 2'h2 == w_state; // @[Mux.scala 80:60]
  wire  _T_22 = 2'h3 == w_state; // @[Mux.scala 80:60]
  wire  isWReq = w_state == 2'h1; // @[AXICache.scala 99:24]
  wire  isWData = w_state == 2'h2; // @[AXICache.scala 100:25]
  wire  isWB = w_state == 2'h3; // @[AXICache.scala 101:22]
  wire  _T_27 = isWReq | isWData; // @[AXICache.scala 126:29]
  assign io_axiIO_awvalid = w_state == 2'h1; // @[AXICache.scala 117:20]
  assign io_axiIO_awaddr = isWReq ? io_cache_w_addr_o : 32'h0; // @[AXICache.scala 118:19]
  assign io_axiIO_awsize = {{1'd0}, io_cache_wsize}; // @[AXICache.scala 121:19]
  assign io_axiIO_wvalid = isWReq | isWData; // @[AXICache.scala 126:19]
  assign io_axiIO_wdata = _T_27 ? io_cache_w_data_o : 64'h0; // @[AXICache.scala 127:18]
  assign io_axiIO_wstrb = _T_27 ? io_cache_w_mask_o : 8'h0; // @[AXICache.scala 128:18]
  assign io_axiIO_wlast = isWReq | isWData; // @[AXICache.scala 129:18]
  assign io_axiIO_bready = w_state == 2'h3; // @[AXICache.scala 132:19]
  assign io_axiIO_arvalid = rd_state == 2'h1; // @[AXICache.scala 58:19]
  assign io_axiIO_araddr = isReq ? io_cache_ar_addr_o : 32'h0; // @[AXICache.scala 59:19]
  assign io_axiIO_arlen = isReq ? io_cache_ar_len_o : 8'h0; // @[AXICache.scala 61:18]
  assign io_axiIO_arsize = {{1'd0}, _T_12}; // @[AXICache.scala 62:19]
  assign io_axiIO_arburst = isReq ? 2'h1 : 2'h0; // @[AXICache.scala 63:20]
  assign io_axiIO_rready = isData | isReq; // @[AXICache.scala 66:18]
  assign io_cache_r_valid_i = io_axiIO_rvalid; // @[AXICache.scala 51:22]
  assign io_cache_r_data_i = io_axiIO_rdata; // @[AXICache.scala 52:21]
  assign io_cache_r_last_i = io_axiIO_rlast; // @[AXICache.scala 50:21]
  assign io_cache_w_ready_i = io_axiIO_bvalid & isWB; // @[AXICache.scala 103:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      rd_state <= 2'h0;
    end else if (_T_7) begin
      if (_T) begin
        rd_state <= 2'h0;
      end else begin
        rd_state <= 2'h2;
      end
    end else if (_T_5) begin
      if (io_axiIO_arready) begin
        if (_T) begin
          rd_state <= 2'h0;
        end else begin
          rd_state <= 2'h2;
        end
      end else begin
        rd_state <= 2'h1;
      end
    end else if (_T_3) begin
      if (io_cache_ar_valid_o) begin
        rd_state <= 2'h1;
      end else begin
        rd_state <= 2'h0;
      end
    end
    if (reset) begin
      w_state <= 2'h0;
    end else if (_T_22) begin
      if (io_axiIO_bvalid) begin
        w_state <= 2'h0;
      end else begin
        w_state <= 2'h3;
      end
    end else if (_T_20) begin
      if (io_axiIO_wready) begin
        w_state <= 2'h3;
      end else begin
        w_state <= 2'h2;
      end
    end else if (_T_18) begin
      if (_T_17) begin
        w_state <= 2'h3;
      end else if (_T_15) begin
        w_state <= 2'h2;
      end else begin
        w_state <= 2'h1;
      end
    end else if (io_cache_w_valid_o) begin
      w_state <= 2'h1;
    end else begin
      w_state <= 2'h0;
    end
  end
endmodule
module arbCpu2DCache(
  input         io_arbIn_valid,
  output        io_arbIn_ready,
  output [63:0] io_arbIn_data_read,
  input  [63:0] io_arbIn_data_write,
  input         io_arbIn_wen,
  input  [31:0] io_arbIn_addr,
  input  [1:0]  io_arbIn_rsize,
  input  [7:0]  io_arbIn_mask,
  output        io_arbMMIO_valid,
  input         io_arbMMIO_ready,
  input  [63:0] io_arbMMIO_data_read,
  output [63:0] io_arbMMIO_data_write,
  output        io_arbMMIO_wen,
  output [31:0] io_arbMMIO_addr,
  output [1:0]  io_arbMMIO_rsize,
  output [7:0]  io_arbMMIO_mask,
  output        io_arbClint_valid,
  input  [63:0] io_arbClint_data_read,
  output [63:0] io_arbClint_data_write,
  output        io_arbClint_wen,
  output [31:0] io_arbClint_addr,
  output        io_arbDCache_valid,
  input         io_arbDCache_ready,
  input  [63:0] io_arbDCache_data_read,
  output [63:0] io_arbDCache_data_write,
  output        io_arbDCache_wen,
  output [31:0] io_arbDCache_addr,
  output [1:0]  io_arbDCache_rsize,
  output [7:0]  io_arbDCache_mask
);
  wire  _T = io_arbIn_addr >= 32'h2000000; // @[arbCpu2Cache.scala 42:31]
  wire  _T_1 = io_arbIn_addr < 32'h200bfff; // @[arbCpu2Cache.scala 42:61]
  wire  clinitV = _T & _T_1; // @[arbCpu2Cache.scala 42:45]
  wire  _T_2 = io_arbIn_addr >= 32'h80000000; // @[arbCpu2Cache.scala 43:31]
  wire  _T_3 = io_arbIn_addr < 32'h8fffffff; // @[arbCpu2Cache.scala 43:60]
  wire  dCacheV = _T_2 & _T_3; // @[arbCpu2Cache.scala 43:44]
  wire  _T_6 = ~clinitV; // @[arbCpu2Cache.scala 47:23]
  wire  _T_7 = ~dCacheV; // @[arbCpu2Cache.scala 47:35]
  wire  _T_8 = _T_6 & _T_7; // @[arbCpu2Cache.scala 47:32]
  wire  _T_11 = dCacheV & io_arbDCache_ready; // @[arbCpu2Cache.scala 56:63]
  wire  _T_12 = clinitV | _T_11; // @[arbCpu2Cache.scala 56:51]
  wire  _T_16 = _T_8 & io_arbMMIO_ready; // @[arbCpu2Cache.scala 56:110]
  wire [63:0] _T_18 = clinitV ? io_arbClint_data_read : io_arbMMIO_data_read; // @[arbCpu2Cache.scala 57:63]
  assign io_arbIn_ready = _T_12 | _T_16; // @[arbCpu2Cache.scala 56:18]
  assign io_arbIn_data_read = dCacheV ? io_arbDCache_data_read : _T_18; // @[arbCpu2Cache.scala 57:22]
  assign io_arbMMIO_valid = _T_8 & io_arbIn_valid; // @[arbCpu2Cache.scala 47:20]
  assign io_arbMMIO_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 50:23]
  assign io_arbClint_valid = clinitV & io_arbIn_valid; // @[arbCpu2Cache.scala 45:21]
  assign io_arbClint_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 51:24]
  assign io_arbClint_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 51:24]
  assign io_arbClint_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 51:24]
  assign io_arbDCache_valid = dCacheV & io_arbIn_valid; // @[arbCpu2Cache.scala 46:22]
  assign io_arbDCache_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 52:25]
endmodule
module mmioCache(
  input         clock,
  input         reset,
  input         io_block,
  input         io_mmioIn_valid,
  output        io_mmioIn_ready,
  output [63:0] io_mmioIn_data_read,
  input  [63:0] io_mmioIn_data_write,
  input         io_mmioIn_wen,
  input  [31:0] io_mmioIn_addr,
  input  [1:0]  io_mmioIn_rsize,
  input  [7:0]  io_mmioIn_mask,
  output        io_mmioOut_valid,
  input         io_mmioOut_ready,
  input  [63:0] io_mmioOut_data_read,
  output [63:0] io_mmioOut_data_write,
  output        io_mmioOut_wen,
  output [31:0] io_mmioOut_addr,
  output [1:0]  io_mmioOut_rsize,
  output [7:0]  io_mmioOut_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[mmioCache.scala 17:22]
  wire  _T = 2'h0 == state; // @[Mux.scala 80:60]
  wire  _T_2 = 2'h1 == state; // @[Mux.scala 80:60]
  wire  _T_4 = 2'h2 == state; // @[Mux.scala 80:60]
  wire  isIdle = state == 2'h0; // @[mmioCache.scala 27:22]
  reg [63:0] _T_7; // @[Reg.scala 27:20]
  assign io_mmioIn_ready = state == 2'h2; // @[mmioCache.scala 39:19]
  assign io_mmioIn_data_read = _T_7; // @[mmioCache.scala 38:23]
  assign io_mmioOut_valid = isIdle & io_mmioIn_valid; // @[mmioCache.scala 31:20]
  assign io_mmioOut_data_write = io_mmioIn_data_write; // @[mmioCache.scala 35:25]
  assign io_mmioOut_wen = io_mmioIn_wen; // @[mmioCache.scala 32:18]
  assign io_mmioOut_addr = io_mmioIn_addr; // @[mmioCache.scala 33:19]
  assign io_mmioOut_rsize = io_mmioIn_rsize; // @[mmioCache.scala 36:20]
  assign io_mmioOut_mask = io_mmioIn_mask; // @[mmioCache.scala 34:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  _T_7 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_4) begin
      if (io_block) begin
        state <= 2'h2;
      end else begin
        state <= 2'h0;
      end
    end else if (_T_2) begin
      if (io_mmioOut_ready) begin
        state <= 2'h2;
      end else begin
        state <= 2'h1;
      end
    end else if (_T) begin
      if (io_mmioIn_valid) begin
        state <= 2'h1;
      end else begin
        state <= 2'h0;
      end
    end else begin
      state <= 2'h0;
    end
    if (reset) begin
      _T_7 <= 64'h0;
    end else if (io_mmioOut_ready) begin
      _T_7 <= io_mmioOut_data_read;
    end
  end
endmodule
module Dcache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output         io_cacheOut_w_valid_o,
  input          io_cacheOut_w_ready_i,
  output [63:0]  io_cacheOut_w_data_o,
  output [31:0]  io_cacheOut_w_addr_o,
  output [7:0]   io_cacheOut_w_mask_o,
  output [1:0]   io_cacheOut_wsize,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [63:0]  io_cacheIn_data_write,
  input          io_cacheIn_wen,
  input  [31:0]  io_cacheIn_addr,
  input  [1:0]   io_cacheIn_rsize,
  input  [7:0]   io_cacheIn_mask,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] offset = io_cacheIn_addr[3:0]; // @[Cache.scala 173:31]
  wire [5:0] index = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  wire [21:0] tag = io_cacheIn_addr[31:10]; // @[Cache.scala 175:28]
  reg [1:0] cacheState; // @[Cache.scala 178:27]
  wire  _T = ~io_block; // @[Cache.scala 182:25]
  wire  _T_1 = io_cacheIn_valid & _T; // @[Cache.scala 182:22]
  wire  _T_260 = 6'h3f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_63_0; // @[Reg.scala 27:20]
  wire  _T_258 = 6'h3e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_62_0; // @[Reg.scala 27:20]
  wire  _T_256 = 6'h3d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_61_0; // @[Reg.scala 27:20]
  wire  _T_254 = 6'h3c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_60_0; // @[Reg.scala 27:20]
  wire  _T_252 = 6'h3b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_59_0; // @[Reg.scala 27:20]
  wire  _T_250 = 6'h3a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_58_0; // @[Reg.scala 27:20]
  wire  _T_248 = 6'h39 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_57_0; // @[Reg.scala 27:20]
  wire  _T_246 = 6'h38 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_56_0; // @[Reg.scala 27:20]
  wire  _T_244 = 6'h37 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_55_0; // @[Reg.scala 27:20]
  wire  _T_242 = 6'h36 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_54_0; // @[Reg.scala 27:20]
  wire  _T_240 = 6'h35 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_53_0; // @[Reg.scala 27:20]
  wire  _T_238 = 6'h34 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_52_0; // @[Reg.scala 27:20]
  wire  _T_236 = 6'h33 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_51_0; // @[Reg.scala 27:20]
  wire  _T_234 = 6'h32 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_50_0; // @[Reg.scala 27:20]
  wire  _T_232 = 6'h31 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_49_0; // @[Reg.scala 27:20]
  wire  _T_230 = 6'h30 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_48_0; // @[Reg.scala 27:20]
  wire  _T_228 = 6'h2f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_47_0; // @[Reg.scala 27:20]
  wire  _T_226 = 6'h2e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_46_0; // @[Reg.scala 27:20]
  wire  _T_224 = 6'h2d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_45_0; // @[Reg.scala 27:20]
  wire  _T_222 = 6'h2c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_44_0; // @[Reg.scala 27:20]
  wire  _T_220 = 6'h2b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_43_0; // @[Reg.scala 27:20]
  wire  _T_218 = 6'h2a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_42_0; // @[Reg.scala 27:20]
  wire  _T_216 = 6'h29 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_41_0; // @[Reg.scala 27:20]
  wire  _T_214 = 6'h28 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_40_0; // @[Reg.scala 27:20]
  wire  _T_212 = 6'h27 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_39_0; // @[Reg.scala 27:20]
  wire  _T_210 = 6'h26 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_38_0; // @[Reg.scala 27:20]
  wire  _T_208 = 6'h25 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_37_0; // @[Reg.scala 27:20]
  wire  _T_206 = 6'h24 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_36_0; // @[Reg.scala 27:20]
  wire  _T_204 = 6'h23 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_35_0; // @[Reg.scala 27:20]
  wire  _T_202 = 6'h22 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_34_0; // @[Reg.scala 27:20]
  wire  _T_200 = 6'h21 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_33_0; // @[Reg.scala 27:20]
  wire  _T_198 = 6'h20 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_32_0; // @[Reg.scala 27:20]
  wire  _T_196 = 6'h1f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_31_0; // @[Reg.scala 27:20]
  wire  _T_194 = 6'h1e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_30_0; // @[Reg.scala 27:20]
  wire  _T_192 = 6'h1d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_29_0; // @[Reg.scala 27:20]
  wire  _T_190 = 6'h1c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_28_0; // @[Reg.scala 27:20]
  wire  _T_188 = 6'h1b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_27_0; // @[Reg.scala 27:20]
  wire  _T_186 = 6'h1a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_26_0; // @[Reg.scala 27:20]
  wire  _T_184 = 6'h19 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_25_0; // @[Reg.scala 27:20]
  wire  _T_182 = 6'h18 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_24_0; // @[Reg.scala 27:20]
  wire  _T_180 = 6'h17 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_23_0; // @[Reg.scala 27:20]
  wire  _T_178 = 6'h16 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_22_0; // @[Reg.scala 27:20]
  wire  _T_176 = 6'h15 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_21_0; // @[Reg.scala 27:20]
  wire  _T_174 = 6'h14 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_20_0; // @[Reg.scala 27:20]
  wire  _T_172 = 6'h13 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_19_0; // @[Reg.scala 27:20]
  wire  _T_170 = 6'h12 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_18_0; // @[Reg.scala 27:20]
  wire  _T_168 = 6'h11 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_17_0; // @[Reg.scala 27:20]
  wire  _T_166 = 6'h10 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_16_0; // @[Reg.scala 27:20]
  wire  _T_164 = 6'hf == index; // @[Mux.scala 80:60]
  reg  vArrayWire_15_0; // @[Reg.scala 27:20]
  wire  _T_162 = 6'he == index; // @[Mux.scala 80:60]
  reg  vArrayWire_14_0; // @[Reg.scala 27:20]
  wire  _T_160 = 6'hd == index; // @[Mux.scala 80:60]
  reg  vArrayWire_13_0; // @[Reg.scala 27:20]
  wire  _T_158 = 6'hc == index; // @[Mux.scala 80:60]
  reg  vArrayWire_12_0; // @[Reg.scala 27:20]
  wire  _T_156 = 6'hb == index; // @[Mux.scala 80:60]
  reg  vArrayWire_11_0; // @[Reg.scala 27:20]
  wire  _T_154 = 6'ha == index; // @[Mux.scala 80:60]
  reg  vArrayWire_10_0; // @[Reg.scala 27:20]
  wire  _T_152 = 6'h9 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_9_0; // @[Reg.scala 27:20]
  wire  _T_150 = 6'h8 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_8_0; // @[Reg.scala 27:20]
  wire  _T_148 = 6'h7 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_7_0; // @[Reg.scala 27:20]
  wire  _T_146 = 6'h6 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_6_0; // @[Reg.scala 27:20]
  wire  _T_144 = 6'h5 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_5_0; // @[Reg.scala 27:20]
  wire  _T_142 = 6'h4 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_4_0; // @[Reg.scala 27:20]
  wire  _T_140 = 6'h3 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_3_0; // @[Reg.scala 27:20]
  wire  _T_138 = 6'h2 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_2_0; // @[Reg.scala 27:20]
  wire  _T_136 = 6'h1 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_1_0; // @[Reg.scala 27:20]
  reg  vArrayWire_0_0; // @[Reg.scala 27:20]
  wire  _T_137_0 = _T_136 ? vArrayWire_1_0 : vArrayWire_0_0; // @[Mux.scala 80:57]
  wire  _T_139_0 = _T_138 ? vArrayWire_2_0 : _T_137_0; // @[Mux.scala 80:57]
  wire  _T_141_0 = _T_140 ? vArrayWire_3_0 : _T_139_0; // @[Mux.scala 80:57]
  wire  _T_143_0 = _T_142 ? vArrayWire_4_0 : _T_141_0; // @[Mux.scala 80:57]
  wire  _T_145_0 = _T_144 ? vArrayWire_5_0 : _T_143_0; // @[Mux.scala 80:57]
  wire  _T_147_0 = _T_146 ? vArrayWire_6_0 : _T_145_0; // @[Mux.scala 80:57]
  wire  _T_149_0 = _T_148 ? vArrayWire_7_0 : _T_147_0; // @[Mux.scala 80:57]
  wire  _T_151_0 = _T_150 ? vArrayWire_8_0 : _T_149_0; // @[Mux.scala 80:57]
  wire  _T_153_0 = _T_152 ? vArrayWire_9_0 : _T_151_0; // @[Mux.scala 80:57]
  wire  _T_155_0 = _T_154 ? vArrayWire_10_0 : _T_153_0; // @[Mux.scala 80:57]
  wire  _T_157_0 = _T_156 ? vArrayWire_11_0 : _T_155_0; // @[Mux.scala 80:57]
  wire  _T_159_0 = _T_158 ? vArrayWire_12_0 : _T_157_0; // @[Mux.scala 80:57]
  wire  _T_161_0 = _T_160 ? vArrayWire_13_0 : _T_159_0; // @[Mux.scala 80:57]
  wire  _T_163_0 = _T_162 ? vArrayWire_14_0 : _T_161_0; // @[Mux.scala 80:57]
  wire  _T_165_0 = _T_164 ? vArrayWire_15_0 : _T_163_0; // @[Mux.scala 80:57]
  wire  _T_167_0 = _T_166 ? vArrayWire_16_0 : _T_165_0; // @[Mux.scala 80:57]
  wire  _T_169_0 = _T_168 ? vArrayWire_17_0 : _T_167_0; // @[Mux.scala 80:57]
  wire  _T_171_0 = _T_170 ? vArrayWire_18_0 : _T_169_0; // @[Mux.scala 80:57]
  wire  _T_173_0 = _T_172 ? vArrayWire_19_0 : _T_171_0; // @[Mux.scala 80:57]
  wire  _T_175_0 = _T_174 ? vArrayWire_20_0 : _T_173_0; // @[Mux.scala 80:57]
  wire  _T_177_0 = _T_176 ? vArrayWire_21_0 : _T_175_0; // @[Mux.scala 80:57]
  wire  _T_179_0 = _T_178 ? vArrayWire_22_0 : _T_177_0; // @[Mux.scala 80:57]
  wire  _T_181_0 = _T_180 ? vArrayWire_23_0 : _T_179_0; // @[Mux.scala 80:57]
  wire  _T_183_0 = _T_182 ? vArrayWire_24_0 : _T_181_0; // @[Mux.scala 80:57]
  wire  _T_185_0 = _T_184 ? vArrayWire_25_0 : _T_183_0; // @[Mux.scala 80:57]
  wire  _T_187_0 = _T_186 ? vArrayWire_26_0 : _T_185_0; // @[Mux.scala 80:57]
  wire  _T_189_0 = _T_188 ? vArrayWire_27_0 : _T_187_0; // @[Mux.scala 80:57]
  wire  _T_191_0 = _T_190 ? vArrayWire_28_0 : _T_189_0; // @[Mux.scala 80:57]
  wire  _T_193_0 = _T_192 ? vArrayWire_29_0 : _T_191_0; // @[Mux.scala 80:57]
  wire  _T_195_0 = _T_194 ? vArrayWire_30_0 : _T_193_0; // @[Mux.scala 80:57]
  wire  _T_197_0 = _T_196 ? vArrayWire_31_0 : _T_195_0; // @[Mux.scala 80:57]
  wire  _T_199_0 = _T_198 ? vArrayWire_32_0 : _T_197_0; // @[Mux.scala 80:57]
  wire  _T_201_0 = _T_200 ? vArrayWire_33_0 : _T_199_0; // @[Mux.scala 80:57]
  wire  _T_203_0 = _T_202 ? vArrayWire_34_0 : _T_201_0; // @[Mux.scala 80:57]
  wire  _T_205_0 = _T_204 ? vArrayWire_35_0 : _T_203_0; // @[Mux.scala 80:57]
  wire  _T_207_0 = _T_206 ? vArrayWire_36_0 : _T_205_0; // @[Mux.scala 80:57]
  wire  _T_209_0 = _T_208 ? vArrayWire_37_0 : _T_207_0; // @[Mux.scala 80:57]
  wire  _T_211_0 = _T_210 ? vArrayWire_38_0 : _T_209_0; // @[Mux.scala 80:57]
  wire  _T_213_0 = _T_212 ? vArrayWire_39_0 : _T_211_0; // @[Mux.scala 80:57]
  wire  _T_215_0 = _T_214 ? vArrayWire_40_0 : _T_213_0; // @[Mux.scala 80:57]
  wire  _T_217_0 = _T_216 ? vArrayWire_41_0 : _T_215_0; // @[Mux.scala 80:57]
  wire  _T_219_0 = _T_218 ? vArrayWire_42_0 : _T_217_0; // @[Mux.scala 80:57]
  wire  _T_221_0 = _T_220 ? vArrayWire_43_0 : _T_219_0; // @[Mux.scala 80:57]
  wire  _T_223_0 = _T_222 ? vArrayWire_44_0 : _T_221_0; // @[Mux.scala 80:57]
  wire  _T_225_0 = _T_224 ? vArrayWire_45_0 : _T_223_0; // @[Mux.scala 80:57]
  wire  _T_227_0 = _T_226 ? vArrayWire_46_0 : _T_225_0; // @[Mux.scala 80:57]
  wire  _T_229_0 = _T_228 ? vArrayWire_47_0 : _T_227_0; // @[Mux.scala 80:57]
  wire  _T_231_0 = _T_230 ? vArrayWire_48_0 : _T_229_0; // @[Mux.scala 80:57]
  wire  _T_233_0 = _T_232 ? vArrayWire_49_0 : _T_231_0; // @[Mux.scala 80:57]
  wire  _T_235_0 = _T_234 ? vArrayWire_50_0 : _T_233_0; // @[Mux.scala 80:57]
  wire  _T_237_0 = _T_236 ? vArrayWire_51_0 : _T_235_0; // @[Mux.scala 80:57]
  wire  _T_239_0 = _T_238 ? vArrayWire_52_0 : _T_237_0; // @[Mux.scala 80:57]
  wire  _T_241_0 = _T_240 ? vArrayWire_53_0 : _T_239_0; // @[Mux.scala 80:57]
  wire  _T_243_0 = _T_242 ? vArrayWire_54_0 : _T_241_0; // @[Mux.scala 80:57]
  wire  _T_245_0 = _T_244 ? vArrayWire_55_0 : _T_243_0; // @[Mux.scala 80:57]
  wire  _T_247_0 = _T_246 ? vArrayWire_56_0 : _T_245_0; // @[Mux.scala 80:57]
  wire  _T_249_0 = _T_248 ? vArrayWire_57_0 : _T_247_0; // @[Mux.scala 80:57]
  wire  _T_251_0 = _T_250 ? vArrayWire_58_0 : _T_249_0; // @[Mux.scala 80:57]
  wire  _T_253_0 = _T_252 ? vArrayWire_59_0 : _T_251_0; // @[Mux.scala 80:57]
  wire  _T_255_0 = _T_254 ? vArrayWire_60_0 : _T_253_0; // @[Mux.scala 80:57]
  wire  _T_257_0 = _T_256 ? vArrayWire_61_0 : _T_255_0; // @[Mux.scala 80:57]
  wire  _T_259_0 = _T_258 ? vArrayWire_62_0 : _T_257_0; // @[Mux.scala 80:57]
  wire  vMuxOut_0 = _T_260 ? vArrayWire_63_0 : _T_259_0; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_0; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_0; // @[Reg.scala 27:20]
  wire [21:0] _T_12_0 = _T_136 ? tagArrayWire_1_0 : tagArrayWire_0_0; // @[Mux.scala 80:57]
  wire [21:0] _T_14_0 = _T_138 ? tagArrayWire_2_0 : _T_12_0; // @[Mux.scala 80:57]
  wire [21:0] _T_16_0 = _T_140 ? tagArrayWire_3_0 : _T_14_0; // @[Mux.scala 80:57]
  wire [21:0] _T_18_0 = _T_142 ? tagArrayWire_4_0 : _T_16_0; // @[Mux.scala 80:57]
  wire [21:0] _T_20_0 = _T_144 ? tagArrayWire_5_0 : _T_18_0; // @[Mux.scala 80:57]
  wire [21:0] _T_22_0 = _T_146 ? tagArrayWire_6_0 : _T_20_0; // @[Mux.scala 80:57]
  wire [21:0] _T_24_0 = _T_148 ? tagArrayWire_7_0 : _T_22_0; // @[Mux.scala 80:57]
  wire [21:0] _T_26_0 = _T_150 ? tagArrayWire_8_0 : _T_24_0; // @[Mux.scala 80:57]
  wire [21:0] _T_28_0 = _T_152 ? tagArrayWire_9_0 : _T_26_0; // @[Mux.scala 80:57]
  wire [21:0] _T_30_0 = _T_154 ? tagArrayWire_10_0 : _T_28_0; // @[Mux.scala 80:57]
  wire [21:0] _T_32_0 = _T_156 ? tagArrayWire_11_0 : _T_30_0; // @[Mux.scala 80:57]
  wire [21:0] _T_34_0 = _T_158 ? tagArrayWire_12_0 : _T_32_0; // @[Mux.scala 80:57]
  wire [21:0] _T_36_0 = _T_160 ? tagArrayWire_13_0 : _T_34_0; // @[Mux.scala 80:57]
  wire [21:0] _T_38_0 = _T_162 ? tagArrayWire_14_0 : _T_36_0; // @[Mux.scala 80:57]
  wire [21:0] _T_40_0 = _T_164 ? tagArrayWire_15_0 : _T_38_0; // @[Mux.scala 80:57]
  wire [21:0] _T_42_0 = _T_166 ? tagArrayWire_16_0 : _T_40_0; // @[Mux.scala 80:57]
  wire [21:0] _T_44_0 = _T_168 ? tagArrayWire_17_0 : _T_42_0; // @[Mux.scala 80:57]
  wire [21:0] _T_46_0 = _T_170 ? tagArrayWire_18_0 : _T_44_0; // @[Mux.scala 80:57]
  wire [21:0] _T_48_0 = _T_172 ? tagArrayWire_19_0 : _T_46_0; // @[Mux.scala 80:57]
  wire [21:0] _T_50_0 = _T_174 ? tagArrayWire_20_0 : _T_48_0; // @[Mux.scala 80:57]
  wire [21:0] _T_52_0 = _T_176 ? tagArrayWire_21_0 : _T_50_0; // @[Mux.scala 80:57]
  wire [21:0] _T_54_0 = _T_178 ? tagArrayWire_22_0 : _T_52_0; // @[Mux.scala 80:57]
  wire [21:0] _T_56_0 = _T_180 ? tagArrayWire_23_0 : _T_54_0; // @[Mux.scala 80:57]
  wire [21:0] _T_58_0 = _T_182 ? tagArrayWire_24_0 : _T_56_0; // @[Mux.scala 80:57]
  wire [21:0] _T_60_0 = _T_184 ? tagArrayWire_25_0 : _T_58_0; // @[Mux.scala 80:57]
  wire [21:0] _T_62_0 = _T_186 ? tagArrayWire_26_0 : _T_60_0; // @[Mux.scala 80:57]
  wire [21:0] _T_64_0 = _T_188 ? tagArrayWire_27_0 : _T_62_0; // @[Mux.scala 80:57]
  wire [21:0] _T_66_0 = _T_190 ? tagArrayWire_28_0 : _T_64_0; // @[Mux.scala 80:57]
  wire [21:0] _T_68_0 = _T_192 ? tagArrayWire_29_0 : _T_66_0; // @[Mux.scala 80:57]
  wire [21:0] _T_70_0 = _T_194 ? tagArrayWire_30_0 : _T_68_0; // @[Mux.scala 80:57]
  wire [21:0] _T_72_0 = _T_196 ? tagArrayWire_31_0 : _T_70_0; // @[Mux.scala 80:57]
  wire [21:0] _T_74_0 = _T_198 ? tagArrayWire_32_0 : _T_72_0; // @[Mux.scala 80:57]
  wire [21:0] _T_76_0 = _T_200 ? tagArrayWire_33_0 : _T_74_0; // @[Mux.scala 80:57]
  wire [21:0] _T_78_0 = _T_202 ? tagArrayWire_34_0 : _T_76_0; // @[Mux.scala 80:57]
  wire [21:0] _T_80_0 = _T_204 ? tagArrayWire_35_0 : _T_78_0; // @[Mux.scala 80:57]
  wire [21:0] _T_82_0 = _T_206 ? tagArrayWire_36_0 : _T_80_0; // @[Mux.scala 80:57]
  wire [21:0] _T_84_0 = _T_208 ? tagArrayWire_37_0 : _T_82_0; // @[Mux.scala 80:57]
  wire [21:0] _T_86_0 = _T_210 ? tagArrayWire_38_0 : _T_84_0; // @[Mux.scala 80:57]
  wire [21:0] _T_88_0 = _T_212 ? tagArrayWire_39_0 : _T_86_0; // @[Mux.scala 80:57]
  wire [21:0] _T_90_0 = _T_214 ? tagArrayWire_40_0 : _T_88_0; // @[Mux.scala 80:57]
  wire [21:0] _T_92_0 = _T_216 ? tagArrayWire_41_0 : _T_90_0; // @[Mux.scala 80:57]
  wire [21:0] _T_94_0 = _T_218 ? tagArrayWire_42_0 : _T_92_0; // @[Mux.scala 80:57]
  wire [21:0] _T_96_0 = _T_220 ? tagArrayWire_43_0 : _T_94_0; // @[Mux.scala 80:57]
  wire [21:0] _T_98_0 = _T_222 ? tagArrayWire_44_0 : _T_96_0; // @[Mux.scala 80:57]
  wire [21:0] _T_100_0 = _T_224 ? tagArrayWire_45_0 : _T_98_0; // @[Mux.scala 80:57]
  wire [21:0] _T_102_0 = _T_226 ? tagArrayWire_46_0 : _T_100_0; // @[Mux.scala 80:57]
  wire [21:0] _T_104_0 = _T_228 ? tagArrayWire_47_0 : _T_102_0; // @[Mux.scala 80:57]
  wire [21:0] _T_106_0 = _T_230 ? tagArrayWire_48_0 : _T_104_0; // @[Mux.scala 80:57]
  wire [21:0] _T_108_0 = _T_232 ? tagArrayWire_49_0 : _T_106_0; // @[Mux.scala 80:57]
  wire [21:0] _T_110_0 = _T_234 ? tagArrayWire_50_0 : _T_108_0; // @[Mux.scala 80:57]
  wire [21:0] _T_112_0 = _T_236 ? tagArrayWire_51_0 : _T_110_0; // @[Mux.scala 80:57]
  wire [21:0] _T_114_0 = _T_238 ? tagArrayWire_52_0 : _T_112_0; // @[Mux.scala 80:57]
  wire [21:0] _T_116_0 = _T_240 ? tagArrayWire_53_0 : _T_114_0; // @[Mux.scala 80:57]
  wire [21:0] _T_118_0 = _T_242 ? tagArrayWire_54_0 : _T_116_0; // @[Mux.scala 80:57]
  wire [21:0] _T_120_0 = _T_244 ? tagArrayWire_55_0 : _T_118_0; // @[Mux.scala 80:57]
  wire [21:0] _T_122_0 = _T_246 ? tagArrayWire_56_0 : _T_120_0; // @[Mux.scala 80:57]
  wire [21:0] _T_124_0 = _T_248 ? tagArrayWire_57_0 : _T_122_0; // @[Mux.scala 80:57]
  wire [21:0] _T_126_0 = _T_250 ? tagArrayWire_58_0 : _T_124_0; // @[Mux.scala 80:57]
  wire [21:0] _T_128_0 = _T_252 ? tagArrayWire_59_0 : _T_126_0; // @[Mux.scala 80:57]
  wire [21:0] _T_130_0 = _T_254 ? tagArrayWire_60_0 : _T_128_0; // @[Mux.scala 80:57]
  wire [21:0] _T_132_0 = _T_256 ? tagArrayWire_61_0 : _T_130_0; // @[Mux.scala 80:57]
  wire [21:0] _T_134_0 = _T_258 ? tagArrayWire_62_0 : _T_132_0; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_0 = _T_260 ? tagArrayWire_63_0 : _T_134_0; // @[Mux.scala 80:57]
  wire  _T_261 = tagMuxOut_0 == tag; // @[Cache.scala 243:76]
  wire  hitArray_0 = vMuxOut_0 & _T_261; // @[Cache.scala 243:60]
  reg  vArrayWire_63_1; // @[Reg.scala 27:20]
  reg  vArrayWire_62_1; // @[Reg.scala 27:20]
  reg  vArrayWire_61_1; // @[Reg.scala 27:20]
  reg  vArrayWire_60_1; // @[Reg.scala 27:20]
  reg  vArrayWire_59_1; // @[Reg.scala 27:20]
  reg  vArrayWire_58_1; // @[Reg.scala 27:20]
  reg  vArrayWire_57_1; // @[Reg.scala 27:20]
  reg  vArrayWire_56_1; // @[Reg.scala 27:20]
  reg  vArrayWire_55_1; // @[Reg.scala 27:20]
  reg  vArrayWire_54_1; // @[Reg.scala 27:20]
  reg  vArrayWire_53_1; // @[Reg.scala 27:20]
  reg  vArrayWire_52_1; // @[Reg.scala 27:20]
  reg  vArrayWire_51_1; // @[Reg.scala 27:20]
  reg  vArrayWire_50_1; // @[Reg.scala 27:20]
  reg  vArrayWire_49_1; // @[Reg.scala 27:20]
  reg  vArrayWire_48_1; // @[Reg.scala 27:20]
  reg  vArrayWire_47_1; // @[Reg.scala 27:20]
  reg  vArrayWire_46_1; // @[Reg.scala 27:20]
  reg  vArrayWire_45_1; // @[Reg.scala 27:20]
  reg  vArrayWire_44_1; // @[Reg.scala 27:20]
  reg  vArrayWire_43_1; // @[Reg.scala 27:20]
  reg  vArrayWire_42_1; // @[Reg.scala 27:20]
  reg  vArrayWire_41_1; // @[Reg.scala 27:20]
  reg  vArrayWire_40_1; // @[Reg.scala 27:20]
  reg  vArrayWire_39_1; // @[Reg.scala 27:20]
  reg  vArrayWire_38_1; // @[Reg.scala 27:20]
  reg  vArrayWire_37_1; // @[Reg.scala 27:20]
  reg  vArrayWire_36_1; // @[Reg.scala 27:20]
  reg  vArrayWire_35_1; // @[Reg.scala 27:20]
  reg  vArrayWire_34_1; // @[Reg.scala 27:20]
  reg  vArrayWire_33_1; // @[Reg.scala 27:20]
  reg  vArrayWire_32_1; // @[Reg.scala 27:20]
  reg  vArrayWire_31_1; // @[Reg.scala 27:20]
  reg  vArrayWire_30_1; // @[Reg.scala 27:20]
  reg  vArrayWire_29_1; // @[Reg.scala 27:20]
  reg  vArrayWire_28_1; // @[Reg.scala 27:20]
  reg  vArrayWire_27_1; // @[Reg.scala 27:20]
  reg  vArrayWire_26_1; // @[Reg.scala 27:20]
  reg  vArrayWire_25_1; // @[Reg.scala 27:20]
  reg  vArrayWire_24_1; // @[Reg.scala 27:20]
  reg  vArrayWire_23_1; // @[Reg.scala 27:20]
  reg  vArrayWire_22_1; // @[Reg.scala 27:20]
  reg  vArrayWire_21_1; // @[Reg.scala 27:20]
  reg  vArrayWire_20_1; // @[Reg.scala 27:20]
  reg  vArrayWire_19_1; // @[Reg.scala 27:20]
  reg  vArrayWire_18_1; // @[Reg.scala 27:20]
  reg  vArrayWire_17_1; // @[Reg.scala 27:20]
  reg  vArrayWire_16_1; // @[Reg.scala 27:20]
  reg  vArrayWire_15_1; // @[Reg.scala 27:20]
  reg  vArrayWire_14_1; // @[Reg.scala 27:20]
  reg  vArrayWire_13_1; // @[Reg.scala 27:20]
  reg  vArrayWire_12_1; // @[Reg.scala 27:20]
  reg  vArrayWire_11_1; // @[Reg.scala 27:20]
  reg  vArrayWire_10_1; // @[Reg.scala 27:20]
  reg  vArrayWire_9_1; // @[Reg.scala 27:20]
  reg  vArrayWire_8_1; // @[Reg.scala 27:20]
  reg  vArrayWire_7_1; // @[Reg.scala 27:20]
  reg  vArrayWire_6_1; // @[Reg.scala 27:20]
  reg  vArrayWire_5_1; // @[Reg.scala 27:20]
  reg  vArrayWire_4_1; // @[Reg.scala 27:20]
  reg  vArrayWire_3_1; // @[Reg.scala 27:20]
  reg  vArrayWire_2_1; // @[Reg.scala 27:20]
  reg  vArrayWire_1_1; // @[Reg.scala 27:20]
  reg  vArrayWire_0_1; // @[Reg.scala 27:20]
  wire  _T_137_1 = _T_136 ? vArrayWire_1_1 : vArrayWire_0_1; // @[Mux.scala 80:57]
  wire  _T_139_1 = _T_138 ? vArrayWire_2_1 : _T_137_1; // @[Mux.scala 80:57]
  wire  _T_141_1 = _T_140 ? vArrayWire_3_1 : _T_139_1; // @[Mux.scala 80:57]
  wire  _T_143_1 = _T_142 ? vArrayWire_4_1 : _T_141_1; // @[Mux.scala 80:57]
  wire  _T_145_1 = _T_144 ? vArrayWire_5_1 : _T_143_1; // @[Mux.scala 80:57]
  wire  _T_147_1 = _T_146 ? vArrayWire_6_1 : _T_145_1; // @[Mux.scala 80:57]
  wire  _T_149_1 = _T_148 ? vArrayWire_7_1 : _T_147_1; // @[Mux.scala 80:57]
  wire  _T_151_1 = _T_150 ? vArrayWire_8_1 : _T_149_1; // @[Mux.scala 80:57]
  wire  _T_153_1 = _T_152 ? vArrayWire_9_1 : _T_151_1; // @[Mux.scala 80:57]
  wire  _T_155_1 = _T_154 ? vArrayWire_10_1 : _T_153_1; // @[Mux.scala 80:57]
  wire  _T_157_1 = _T_156 ? vArrayWire_11_1 : _T_155_1; // @[Mux.scala 80:57]
  wire  _T_159_1 = _T_158 ? vArrayWire_12_1 : _T_157_1; // @[Mux.scala 80:57]
  wire  _T_161_1 = _T_160 ? vArrayWire_13_1 : _T_159_1; // @[Mux.scala 80:57]
  wire  _T_163_1 = _T_162 ? vArrayWire_14_1 : _T_161_1; // @[Mux.scala 80:57]
  wire  _T_165_1 = _T_164 ? vArrayWire_15_1 : _T_163_1; // @[Mux.scala 80:57]
  wire  _T_167_1 = _T_166 ? vArrayWire_16_1 : _T_165_1; // @[Mux.scala 80:57]
  wire  _T_169_1 = _T_168 ? vArrayWire_17_1 : _T_167_1; // @[Mux.scala 80:57]
  wire  _T_171_1 = _T_170 ? vArrayWire_18_1 : _T_169_1; // @[Mux.scala 80:57]
  wire  _T_173_1 = _T_172 ? vArrayWire_19_1 : _T_171_1; // @[Mux.scala 80:57]
  wire  _T_175_1 = _T_174 ? vArrayWire_20_1 : _T_173_1; // @[Mux.scala 80:57]
  wire  _T_177_1 = _T_176 ? vArrayWire_21_1 : _T_175_1; // @[Mux.scala 80:57]
  wire  _T_179_1 = _T_178 ? vArrayWire_22_1 : _T_177_1; // @[Mux.scala 80:57]
  wire  _T_181_1 = _T_180 ? vArrayWire_23_1 : _T_179_1; // @[Mux.scala 80:57]
  wire  _T_183_1 = _T_182 ? vArrayWire_24_1 : _T_181_1; // @[Mux.scala 80:57]
  wire  _T_185_1 = _T_184 ? vArrayWire_25_1 : _T_183_1; // @[Mux.scala 80:57]
  wire  _T_187_1 = _T_186 ? vArrayWire_26_1 : _T_185_1; // @[Mux.scala 80:57]
  wire  _T_189_1 = _T_188 ? vArrayWire_27_1 : _T_187_1; // @[Mux.scala 80:57]
  wire  _T_191_1 = _T_190 ? vArrayWire_28_1 : _T_189_1; // @[Mux.scala 80:57]
  wire  _T_193_1 = _T_192 ? vArrayWire_29_1 : _T_191_1; // @[Mux.scala 80:57]
  wire  _T_195_1 = _T_194 ? vArrayWire_30_1 : _T_193_1; // @[Mux.scala 80:57]
  wire  _T_197_1 = _T_196 ? vArrayWire_31_1 : _T_195_1; // @[Mux.scala 80:57]
  wire  _T_199_1 = _T_198 ? vArrayWire_32_1 : _T_197_1; // @[Mux.scala 80:57]
  wire  _T_201_1 = _T_200 ? vArrayWire_33_1 : _T_199_1; // @[Mux.scala 80:57]
  wire  _T_203_1 = _T_202 ? vArrayWire_34_1 : _T_201_1; // @[Mux.scala 80:57]
  wire  _T_205_1 = _T_204 ? vArrayWire_35_1 : _T_203_1; // @[Mux.scala 80:57]
  wire  _T_207_1 = _T_206 ? vArrayWire_36_1 : _T_205_1; // @[Mux.scala 80:57]
  wire  _T_209_1 = _T_208 ? vArrayWire_37_1 : _T_207_1; // @[Mux.scala 80:57]
  wire  _T_211_1 = _T_210 ? vArrayWire_38_1 : _T_209_1; // @[Mux.scala 80:57]
  wire  _T_213_1 = _T_212 ? vArrayWire_39_1 : _T_211_1; // @[Mux.scala 80:57]
  wire  _T_215_1 = _T_214 ? vArrayWire_40_1 : _T_213_1; // @[Mux.scala 80:57]
  wire  _T_217_1 = _T_216 ? vArrayWire_41_1 : _T_215_1; // @[Mux.scala 80:57]
  wire  _T_219_1 = _T_218 ? vArrayWire_42_1 : _T_217_1; // @[Mux.scala 80:57]
  wire  _T_221_1 = _T_220 ? vArrayWire_43_1 : _T_219_1; // @[Mux.scala 80:57]
  wire  _T_223_1 = _T_222 ? vArrayWire_44_1 : _T_221_1; // @[Mux.scala 80:57]
  wire  _T_225_1 = _T_224 ? vArrayWire_45_1 : _T_223_1; // @[Mux.scala 80:57]
  wire  _T_227_1 = _T_226 ? vArrayWire_46_1 : _T_225_1; // @[Mux.scala 80:57]
  wire  _T_229_1 = _T_228 ? vArrayWire_47_1 : _T_227_1; // @[Mux.scala 80:57]
  wire  _T_231_1 = _T_230 ? vArrayWire_48_1 : _T_229_1; // @[Mux.scala 80:57]
  wire  _T_233_1 = _T_232 ? vArrayWire_49_1 : _T_231_1; // @[Mux.scala 80:57]
  wire  _T_235_1 = _T_234 ? vArrayWire_50_1 : _T_233_1; // @[Mux.scala 80:57]
  wire  _T_237_1 = _T_236 ? vArrayWire_51_1 : _T_235_1; // @[Mux.scala 80:57]
  wire  _T_239_1 = _T_238 ? vArrayWire_52_1 : _T_237_1; // @[Mux.scala 80:57]
  wire  _T_241_1 = _T_240 ? vArrayWire_53_1 : _T_239_1; // @[Mux.scala 80:57]
  wire  _T_243_1 = _T_242 ? vArrayWire_54_1 : _T_241_1; // @[Mux.scala 80:57]
  wire  _T_245_1 = _T_244 ? vArrayWire_55_1 : _T_243_1; // @[Mux.scala 80:57]
  wire  _T_247_1 = _T_246 ? vArrayWire_56_1 : _T_245_1; // @[Mux.scala 80:57]
  wire  _T_249_1 = _T_248 ? vArrayWire_57_1 : _T_247_1; // @[Mux.scala 80:57]
  wire  _T_251_1 = _T_250 ? vArrayWire_58_1 : _T_249_1; // @[Mux.scala 80:57]
  wire  _T_253_1 = _T_252 ? vArrayWire_59_1 : _T_251_1; // @[Mux.scala 80:57]
  wire  _T_255_1 = _T_254 ? vArrayWire_60_1 : _T_253_1; // @[Mux.scala 80:57]
  wire  _T_257_1 = _T_256 ? vArrayWire_61_1 : _T_255_1; // @[Mux.scala 80:57]
  wire  _T_259_1 = _T_258 ? vArrayWire_62_1 : _T_257_1; // @[Mux.scala 80:57]
  wire  vMuxOut_1 = _T_260 ? vArrayWire_63_1 : _T_259_1; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_1; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_1; // @[Reg.scala 27:20]
  wire [21:0] _T_12_1 = _T_136 ? tagArrayWire_1_1 : tagArrayWire_0_1; // @[Mux.scala 80:57]
  wire [21:0] _T_14_1 = _T_138 ? tagArrayWire_2_1 : _T_12_1; // @[Mux.scala 80:57]
  wire [21:0] _T_16_1 = _T_140 ? tagArrayWire_3_1 : _T_14_1; // @[Mux.scala 80:57]
  wire [21:0] _T_18_1 = _T_142 ? tagArrayWire_4_1 : _T_16_1; // @[Mux.scala 80:57]
  wire [21:0] _T_20_1 = _T_144 ? tagArrayWire_5_1 : _T_18_1; // @[Mux.scala 80:57]
  wire [21:0] _T_22_1 = _T_146 ? tagArrayWire_6_1 : _T_20_1; // @[Mux.scala 80:57]
  wire [21:0] _T_24_1 = _T_148 ? tagArrayWire_7_1 : _T_22_1; // @[Mux.scala 80:57]
  wire [21:0] _T_26_1 = _T_150 ? tagArrayWire_8_1 : _T_24_1; // @[Mux.scala 80:57]
  wire [21:0] _T_28_1 = _T_152 ? tagArrayWire_9_1 : _T_26_1; // @[Mux.scala 80:57]
  wire [21:0] _T_30_1 = _T_154 ? tagArrayWire_10_1 : _T_28_1; // @[Mux.scala 80:57]
  wire [21:0] _T_32_1 = _T_156 ? tagArrayWire_11_1 : _T_30_1; // @[Mux.scala 80:57]
  wire [21:0] _T_34_1 = _T_158 ? tagArrayWire_12_1 : _T_32_1; // @[Mux.scala 80:57]
  wire [21:0] _T_36_1 = _T_160 ? tagArrayWire_13_1 : _T_34_1; // @[Mux.scala 80:57]
  wire [21:0] _T_38_1 = _T_162 ? tagArrayWire_14_1 : _T_36_1; // @[Mux.scala 80:57]
  wire [21:0] _T_40_1 = _T_164 ? tagArrayWire_15_1 : _T_38_1; // @[Mux.scala 80:57]
  wire [21:0] _T_42_1 = _T_166 ? tagArrayWire_16_1 : _T_40_1; // @[Mux.scala 80:57]
  wire [21:0] _T_44_1 = _T_168 ? tagArrayWire_17_1 : _T_42_1; // @[Mux.scala 80:57]
  wire [21:0] _T_46_1 = _T_170 ? tagArrayWire_18_1 : _T_44_1; // @[Mux.scala 80:57]
  wire [21:0] _T_48_1 = _T_172 ? tagArrayWire_19_1 : _T_46_1; // @[Mux.scala 80:57]
  wire [21:0] _T_50_1 = _T_174 ? tagArrayWire_20_1 : _T_48_1; // @[Mux.scala 80:57]
  wire [21:0] _T_52_1 = _T_176 ? tagArrayWire_21_1 : _T_50_1; // @[Mux.scala 80:57]
  wire [21:0] _T_54_1 = _T_178 ? tagArrayWire_22_1 : _T_52_1; // @[Mux.scala 80:57]
  wire [21:0] _T_56_1 = _T_180 ? tagArrayWire_23_1 : _T_54_1; // @[Mux.scala 80:57]
  wire [21:0] _T_58_1 = _T_182 ? tagArrayWire_24_1 : _T_56_1; // @[Mux.scala 80:57]
  wire [21:0] _T_60_1 = _T_184 ? tagArrayWire_25_1 : _T_58_1; // @[Mux.scala 80:57]
  wire [21:0] _T_62_1 = _T_186 ? tagArrayWire_26_1 : _T_60_1; // @[Mux.scala 80:57]
  wire [21:0] _T_64_1 = _T_188 ? tagArrayWire_27_1 : _T_62_1; // @[Mux.scala 80:57]
  wire [21:0] _T_66_1 = _T_190 ? tagArrayWire_28_1 : _T_64_1; // @[Mux.scala 80:57]
  wire [21:0] _T_68_1 = _T_192 ? tagArrayWire_29_1 : _T_66_1; // @[Mux.scala 80:57]
  wire [21:0] _T_70_1 = _T_194 ? tagArrayWire_30_1 : _T_68_1; // @[Mux.scala 80:57]
  wire [21:0] _T_72_1 = _T_196 ? tagArrayWire_31_1 : _T_70_1; // @[Mux.scala 80:57]
  wire [21:0] _T_74_1 = _T_198 ? tagArrayWire_32_1 : _T_72_1; // @[Mux.scala 80:57]
  wire [21:0] _T_76_1 = _T_200 ? tagArrayWire_33_1 : _T_74_1; // @[Mux.scala 80:57]
  wire [21:0] _T_78_1 = _T_202 ? tagArrayWire_34_1 : _T_76_1; // @[Mux.scala 80:57]
  wire [21:0] _T_80_1 = _T_204 ? tagArrayWire_35_1 : _T_78_1; // @[Mux.scala 80:57]
  wire [21:0] _T_82_1 = _T_206 ? tagArrayWire_36_1 : _T_80_1; // @[Mux.scala 80:57]
  wire [21:0] _T_84_1 = _T_208 ? tagArrayWire_37_1 : _T_82_1; // @[Mux.scala 80:57]
  wire [21:0] _T_86_1 = _T_210 ? tagArrayWire_38_1 : _T_84_1; // @[Mux.scala 80:57]
  wire [21:0] _T_88_1 = _T_212 ? tagArrayWire_39_1 : _T_86_1; // @[Mux.scala 80:57]
  wire [21:0] _T_90_1 = _T_214 ? tagArrayWire_40_1 : _T_88_1; // @[Mux.scala 80:57]
  wire [21:0] _T_92_1 = _T_216 ? tagArrayWire_41_1 : _T_90_1; // @[Mux.scala 80:57]
  wire [21:0] _T_94_1 = _T_218 ? tagArrayWire_42_1 : _T_92_1; // @[Mux.scala 80:57]
  wire [21:0] _T_96_1 = _T_220 ? tagArrayWire_43_1 : _T_94_1; // @[Mux.scala 80:57]
  wire [21:0] _T_98_1 = _T_222 ? tagArrayWire_44_1 : _T_96_1; // @[Mux.scala 80:57]
  wire [21:0] _T_100_1 = _T_224 ? tagArrayWire_45_1 : _T_98_1; // @[Mux.scala 80:57]
  wire [21:0] _T_102_1 = _T_226 ? tagArrayWire_46_1 : _T_100_1; // @[Mux.scala 80:57]
  wire [21:0] _T_104_1 = _T_228 ? tagArrayWire_47_1 : _T_102_1; // @[Mux.scala 80:57]
  wire [21:0] _T_106_1 = _T_230 ? tagArrayWire_48_1 : _T_104_1; // @[Mux.scala 80:57]
  wire [21:0] _T_108_1 = _T_232 ? tagArrayWire_49_1 : _T_106_1; // @[Mux.scala 80:57]
  wire [21:0] _T_110_1 = _T_234 ? tagArrayWire_50_1 : _T_108_1; // @[Mux.scala 80:57]
  wire [21:0] _T_112_1 = _T_236 ? tagArrayWire_51_1 : _T_110_1; // @[Mux.scala 80:57]
  wire [21:0] _T_114_1 = _T_238 ? tagArrayWire_52_1 : _T_112_1; // @[Mux.scala 80:57]
  wire [21:0] _T_116_1 = _T_240 ? tagArrayWire_53_1 : _T_114_1; // @[Mux.scala 80:57]
  wire [21:0] _T_118_1 = _T_242 ? tagArrayWire_54_1 : _T_116_1; // @[Mux.scala 80:57]
  wire [21:0] _T_120_1 = _T_244 ? tagArrayWire_55_1 : _T_118_1; // @[Mux.scala 80:57]
  wire [21:0] _T_122_1 = _T_246 ? tagArrayWire_56_1 : _T_120_1; // @[Mux.scala 80:57]
  wire [21:0] _T_124_1 = _T_248 ? tagArrayWire_57_1 : _T_122_1; // @[Mux.scala 80:57]
  wire [21:0] _T_126_1 = _T_250 ? tagArrayWire_58_1 : _T_124_1; // @[Mux.scala 80:57]
  wire [21:0] _T_128_1 = _T_252 ? tagArrayWire_59_1 : _T_126_1; // @[Mux.scala 80:57]
  wire [21:0] _T_130_1 = _T_254 ? tagArrayWire_60_1 : _T_128_1; // @[Mux.scala 80:57]
  wire [21:0] _T_132_1 = _T_256 ? tagArrayWire_61_1 : _T_130_1; // @[Mux.scala 80:57]
  wire [21:0] _T_134_1 = _T_258 ? tagArrayWire_62_1 : _T_132_1; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_1 = _T_260 ? tagArrayWire_63_1 : _T_134_1; // @[Mux.scala 80:57]
  wire  _T_262 = tagMuxOut_1 == tag; // @[Cache.scala 243:76]
  wire  hitArray_1 = vMuxOut_1 & _T_262; // @[Cache.scala 243:60]
  wire  _T_266 = hitArray_0 | hitArray_1; // @[Cache.scala 244:49]
  reg  vArrayWire_63_2; // @[Reg.scala 27:20]
  reg  vArrayWire_62_2; // @[Reg.scala 27:20]
  reg  vArrayWire_61_2; // @[Reg.scala 27:20]
  reg  vArrayWire_60_2; // @[Reg.scala 27:20]
  reg  vArrayWire_59_2; // @[Reg.scala 27:20]
  reg  vArrayWire_58_2; // @[Reg.scala 27:20]
  reg  vArrayWire_57_2; // @[Reg.scala 27:20]
  reg  vArrayWire_56_2; // @[Reg.scala 27:20]
  reg  vArrayWire_55_2; // @[Reg.scala 27:20]
  reg  vArrayWire_54_2; // @[Reg.scala 27:20]
  reg  vArrayWire_53_2; // @[Reg.scala 27:20]
  reg  vArrayWire_52_2; // @[Reg.scala 27:20]
  reg  vArrayWire_51_2; // @[Reg.scala 27:20]
  reg  vArrayWire_50_2; // @[Reg.scala 27:20]
  reg  vArrayWire_49_2; // @[Reg.scala 27:20]
  reg  vArrayWire_48_2; // @[Reg.scala 27:20]
  reg  vArrayWire_47_2; // @[Reg.scala 27:20]
  reg  vArrayWire_46_2; // @[Reg.scala 27:20]
  reg  vArrayWire_45_2; // @[Reg.scala 27:20]
  reg  vArrayWire_44_2; // @[Reg.scala 27:20]
  reg  vArrayWire_43_2; // @[Reg.scala 27:20]
  reg  vArrayWire_42_2; // @[Reg.scala 27:20]
  reg  vArrayWire_41_2; // @[Reg.scala 27:20]
  reg  vArrayWire_40_2; // @[Reg.scala 27:20]
  reg  vArrayWire_39_2; // @[Reg.scala 27:20]
  reg  vArrayWire_38_2; // @[Reg.scala 27:20]
  reg  vArrayWire_37_2; // @[Reg.scala 27:20]
  reg  vArrayWire_36_2; // @[Reg.scala 27:20]
  reg  vArrayWire_35_2; // @[Reg.scala 27:20]
  reg  vArrayWire_34_2; // @[Reg.scala 27:20]
  reg  vArrayWire_33_2; // @[Reg.scala 27:20]
  reg  vArrayWire_32_2; // @[Reg.scala 27:20]
  reg  vArrayWire_31_2; // @[Reg.scala 27:20]
  reg  vArrayWire_30_2; // @[Reg.scala 27:20]
  reg  vArrayWire_29_2; // @[Reg.scala 27:20]
  reg  vArrayWire_28_2; // @[Reg.scala 27:20]
  reg  vArrayWire_27_2; // @[Reg.scala 27:20]
  reg  vArrayWire_26_2; // @[Reg.scala 27:20]
  reg  vArrayWire_25_2; // @[Reg.scala 27:20]
  reg  vArrayWire_24_2; // @[Reg.scala 27:20]
  reg  vArrayWire_23_2; // @[Reg.scala 27:20]
  reg  vArrayWire_22_2; // @[Reg.scala 27:20]
  reg  vArrayWire_21_2; // @[Reg.scala 27:20]
  reg  vArrayWire_20_2; // @[Reg.scala 27:20]
  reg  vArrayWire_19_2; // @[Reg.scala 27:20]
  reg  vArrayWire_18_2; // @[Reg.scala 27:20]
  reg  vArrayWire_17_2; // @[Reg.scala 27:20]
  reg  vArrayWire_16_2; // @[Reg.scala 27:20]
  reg  vArrayWire_15_2; // @[Reg.scala 27:20]
  reg  vArrayWire_14_2; // @[Reg.scala 27:20]
  reg  vArrayWire_13_2; // @[Reg.scala 27:20]
  reg  vArrayWire_12_2; // @[Reg.scala 27:20]
  reg  vArrayWire_11_2; // @[Reg.scala 27:20]
  reg  vArrayWire_10_2; // @[Reg.scala 27:20]
  reg  vArrayWire_9_2; // @[Reg.scala 27:20]
  reg  vArrayWire_8_2; // @[Reg.scala 27:20]
  reg  vArrayWire_7_2; // @[Reg.scala 27:20]
  reg  vArrayWire_6_2; // @[Reg.scala 27:20]
  reg  vArrayWire_5_2; // @[Reg.scala 27:20]
  reg  vArrayWire_4_2; // @[Reg.scala 27:20]
  reg  vArrayWire_3_2; // @[Reg.scala 27:20]
  reg  vArrayWire_2_2; // @[Reg.scala 27:20]
  reg  vArrayWire_1_2; // @[Reg.scala 27:20]
  reg  vArrayWire_0_2; // @[Reg.scala 27:20]
  wire  _T_137_2 = _T_136 ? vArrayWire_1_2 : vArrayWire_0_2; // @[Mux.scala 80:57]
  wire  _T_139_2 = _T_138 ? vArrayWire_2_2 : _T_137_2; // @[Mux.scala 80:57]
  wire  _T_141_2 = _T_140 ? vArrayWire_3_2 : _T_139_2; // @[Mux.scala 80:57]
  wire  _T_143_2 = _T_142 ? vArrayWire_4_2 : _T_141_2; // @[Mux.scala 80:57]
  wire  _T_145_2 = _T_144 ? vArrayWire_5_2 : _T_143_2; // @[Mux.scala 80:57]
  wire  _T_147_2 = _T_146 ? vArrayWire_6_2 : _T_145_2; // @[Mux.scala 80:57]
  wire  _T_149_2 = _T_148 ? vArrayWire_7_2 : _T_147_2; // @[Mux.scala 80:57]
  wire  _T_151_2 = _T_150 ? vArrayWire_8_2 : _T_149_2; // @[Mux.scala 80:57]
  wire  _T_153_2 = _T_152 ? vArrayWire_9_2 : _T_151_2; // @[Mux.scala 80:57]
  wire  _T_155_2 = _T_154 ? vArrayWire_10_2 : _T_153_2; // @[Mux.scala 80:57]
  wire  _T_157_2 = _T_156 ? vArrayWire_11_2 : _T_155_2; // @[Mux.scala 80:57]
  wire  _T_159_2 = _T_158 ? vArrayWire_12_2 : _T_157_2; // @[Mux.scala 80:57]
  wire  _T_161_2 = _T_160 ? vArrayWire_13_2 : _T_159_2; // @[Mux.scala 80:57]
  wire  _T_163_2 = _T_162 ? vArrayWire_14_2 : _T_161_2; // @[Mux.scala 80:57]
  wire  _T_165_2 = _T_164 ? vArrayWire_15_2 : _T_163_2; // @[Mux.scala 80:57]
  wire  _T_167_2 = _T_166 ? vArrayWire_16_2 : _T_165_2; // @[Mux.scala 80:57]
  wire  _T_169_2 = _T_168 ? vArrayWire_17_2 : _T_167_2; // @[Mux.scala 80:57]
  wire  _T_171_2 = _T_170 ? vArrayWire_18_2 : _T_169_2; // @[Mux.scala 80:57]
  wire  _T_173_2 = _T_172 ? vArrayWire_19_2 : _T_171_2; // @[Mux.scala 80:57]
  wire  _T_175_2 = _T_174 ? vArrayWire_20_2 : _T_173_2; // @[Mux.scala 80:57]
  wire  _T_177_2 = _T_176 ? vArrayWire_21_2 : _T_175_2; // @[Mux.scala 80:57]
  wire  _T_179_2 = _T_178 ? vArrayWire_22_2 : _T_177_2; // @[Mux.scala 80:57]
  wire  _T_181_2 = _T_180 ? vArrayWire_23_2 : _T_179_2; // @[Mux.scala 80:57]
  wire  _T_183_2 = _T_182 ? vArrayWire_24_2 : _T_181_2; // @[Mux.scala 80:57]
  wire  _T_185_2 = _T_184 ? vArrayWire_25_2 : _T_183_2; // @[Mux.scala 80:57]
  wire  _T_187_2 = _T_186 ? vArrayWire_26_2 : _T_185_2; // @[Mux.scala 80:57]
  wire  _T_189_2 = _T_188 ? vArrayWire_27_2 : _T_187_2; // @[Mux.scala 80:57]
  wire  _T_191_2 = _T_190 ? vArrayWire_28_2 : _T_189_2; // @[Mux.scala 80:57]
  wire  _T_193_2 = _T_192 ? vArrayWire_29_2 : _T_191_2; // @[Mux.scala 80:57]
  wire  _T_195_2 = _T_194 ? vArrayWire_30_2 : _T_193_2; // @[Mux.scala 80:57]
  wire  _T_197_2 = _T_196 ? vArrayWire_31_2 : _T_195_2; // @[Mux.scala 80:57]
  wire  _T_199_2 = _T_198 ? vArrayWire_32_2 : _T_197_2; // @[Mux.scala 80:57]
  wire  _T_201_2 = _T_200 ? vArrayWire_33_2 : _T_199_2; // @[Mux.scala 80:57]
  wire  _T_203_2 = _T_202 ? vArrayWire_34_2 : _T_201_2; // @[Mux.scala 80:57]
  wire  _T_205_2 = _T_204 ? vArrayWire_35_2 : _T_203_2; // @[Mux.scala 80:57]
  wire  _T_207_2 = _T_206 ? vArrayWire_36_2 : _T_205_2; // @[Mux.scala 80:57]
  wire  _T_209_2 = _T_208 ? vArrayWire_37_2 : _T_207_2; // @[Mux.scala 80:57]
  wire  _T_211_2 = _T_210 ? vArrayWire_38_2 : _T_209_2; // @[Mux.scala 80:57]
  wire  _T_213_2 = _T_212 ? vArrayWire_39_2 : _T_211_2; // @[Mux.scala 80:57]
  wire  _T_215_2 = _T_214 ? vArrayWire_40_2 : _T_213_2; // @[Mux.scala 80:57]
  wire  _T_217_2 = _T_216 ? vArrayWire_41_2 : _T_215_2; // @[Mux.scala 80:57]
  wire  _T_219_2 = _T_218 ? vArrayWire_42_2 : _T_217_2; // @[Mux.scala 80:57]
  wire  _T_221_2 = _T_220 ? vArrayWire_43_2 : _T_219_2; // @[Mux.scala 80:57]
  wire  _T_223_2 = _T_222 ? vArrayWire_44_2 : _T_221_2; // @[Mux.scala 80:57]
  wire  _T_225_2 = _T_224 ? vArrayWire_45_2 : _T_223_2; // @[Mux.scala 80:57]
  wire  _T_227_2 = _T_226 ? vArrayWire_46_2 : _T_225_2; // @[Mux.scala 80:57]
  wire  _T_229_2 = _T_228 ? vArrayWire_47_2 : _T_227_2; // @[Mux.scala 80:57]
  wire  _T_231_2 = _T_230 ? vArrayWire_48_2 : _T_229_2; // @[Mux.scala 80:57]
  wire  _T_233_2 = _T_232 ? vArrayWire_49_2 : _T_231_2; // @[Mux.scala 80:57]
  wire  _T_235_2 = _T_234 ? vArrayWire_50_2 : _T_233_2; // @[Mux.scala 80:57]
  wire  _T_237_2 = _T_236 ? vArrayWire_51_2 : _T_235_2; // @[Mux.scala 80:57]
  wire  _T_239_2 = _T_238 ? vArrayWire_52_2 : _T_237_2; // @[Mux.scala 80:57]
  wire  _T_241_2 = _T_240 ? vArrayWire_53_2 : _T_239_2; // @[Mux.scala 80:57]
  wire  _T_243_2 = _T_242 ? vArrayWire_54_2 : _T_241_2; // @[Mux.scala 80:57]
  wire  _T_245_2 = _T_244 ? vArrayWire_55_2 : _T_243_2; // @[Mux.scala 80:57]
  wire  _T_247_2 = _T_246 ? vArrayWire_56_2 : _T_245_2; // @[Mux.scala 80:57]
  wire  _T_249_2 = _T_248 ? vArrayWire_57_2 : _T_247_2; // @[Mux.scala 80:57]
  wire  _T_251_2 = _T_250 ? vArrayWire_58_2 : _T_249_2; // @[Mux.scala 80:57]
  wire  _T_253_2 = _T_252 ? vArrayWire_59_2 : _T_251_2; // @[Mux.scala 80:57]
  wire  _T_255_2 = _T_254 ? vArrayWire_60_2 : _T_253_2; // @[Mux.scala 80:57]
  wire  _T_257_2 = _T_256 ? vArrayWire_61_2 : _T_255_2; // @[Mux.scala 80:57]
  wire  _T_259_2 = _T_258 ? vArrayWire_62_2 : _T_257_2; // @[Mux.scala 80:57]
  wire  vMuxOut_2 = _T_260 ? vArrayWire_63_2 : _T_259_2; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_2; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_2; // @[Reg.scala 27:20]
  wire [21:0] _T_12_2 = _T_136 ? tagArrayWire_1_2 : tagArrayWire_0_2; // @[Mux.scala 80:57]
  wire [21:0] _T_14_2 = _T_138 ? tagArrayWire_2_2 : _T_12_2; // @[Mux.scala 80:57]
  wire [21:0] _T_16_2 = _T_140 ? tagArrayWire_3_2 : _T_14_2; // @[Mux.scala 80:57]
  wire [21:0] _T_18_2 = _T_142 ? tagArrayWire_4_2 : _T_16_2; // @[Mux.scala 80:57]
  wire [21:0] _T_20_2 = _T_144 ? tagArrayWire_5_2 : _T_18_2; // @[Mux.scala 80:57]
  wire [21:0] _T_22_2 = _T_146 ? tagArrayWire_6_2 : _T_20_2; // @[Mux.scala 80:57]
  wire [21:0] _T_24_2 = _T_148 ? tagArrayWire_7_2 : _T_22_2; // @[Mux.scala 80:57]
  wire [21:0] _T_26_2 = _T_150 ? tagArrayWire_8_2 : _T_24_2; // @[Mux.scala 80:57]
  wire [21:0] _T_28_2 = _T_152 ? tagArrayWire_9_2 : _T_26_2; // @[Mux.scala 80:57]
  wire [21:0] _T_30_2 = _T_154 ? tagArrayWire_10_2 : _T_28_2; // @[Mux.scala 80:57]
  wire [21:0] _T_32_2 = _T_156 ? tagArrayWire_11_2 : _T_30_2; // @[Mux.scala 80:57]
  wire [21:0] _T_34_2 = _T_158 ? tagArrayWire_12_2 : _T_32_2; // @[Mux.scala 80:57]
  wire [21:0] _T_36_2 = _T_160 ? tagArrayWire_13_2 : _T_34_2; // @[Mux.scala 80:57]
  wire [21:0] _T_38_2 = _T_162 ? tagArrayWire_14_2 : _T_36_2; // @[Mux.scala 80:57]
  wire [21:0] _T_40_2 = _T_164 ? tagArrayWire_15_2 : _T_38_2; // @[Mux.scala 80:57]
  wire [21:0] _T_42_2 = _T_166 ? tagArrayWire_16_2 : _T_40_2; // @[Mux.scala 80:57]
  wire [21:0] _T_44_2 = _T_168 ? tagArrayWire_17_2 : _T_42_2; // @[Mux.scala 80:57]
  wire [21:0] _T_46_2 = _T_170 ? tagArrayWire_18_2 : _T_44_2; // @[Mux.scala 80:57]
  wire [21:0] _T_48_2 = _T_172 ? tagArrayWire_19_2 : _T_46_2; // @[Mux.scala 80:57]
  wire [21:0] _T_50_2 = _T_174 ? tagArrayWire_20_2 : _T_48_2; // @[Mux.scala 80:57]
  wire [21:0] _T_52_2 = _T_176 ? tagArrayWire_21_2 : _T_50_2; // @[Mux.scala 80:57]
  wire [21:0] _T_54_2 = _T_178 ? tagArrayWire_22_2 : _T_52_2; // @[Mux.scala 80:57]
  wire [21:0] _T_56_2 = _T_180 ? tagArrayWire_23_2 : _T_54_2; // @[Mux.scala 80:57]
  wire [21:0] _T_58_2 = _T_182 ? tagArrayWire_24_2 : _T_56_2; // @[Mux.scala 80:57]
  wire [21:0] _T_60_2 = _T_184 ? tagArrayWire_25_2 : _T_58_2; // @[Mux.scala 80:57]
  wire [21:0] _T_62_2 = _T_186 ? tagArrayWire_26_2 : _T_60_2; // @[Mux.scala 80:57]
  wire [21:0] _T_64_2 = _T_188 ? tagArrayWire_27_2 : _T_62_2; // @[Mux.scala 80:57]
  wire [21:0] _T_66_2 = _T_190 ? tagArrayWire_28_2 : _T_64_2; // @[Mux.scala 80:57]
  wire [21:0] _T_68_2 = _T_192 ? tagArrayWire_29_2 : _T_66_2; // @[Mux.scala 80:57]
  wire [21:0] _T_70_2 = _T_194 ? tagArrayWire_30_2 : _T_68_2; // @[Mux.scala 80:57]
  wire [21:0] _T_72_2 = _T_196 ? tagArrayWire_31_2 : _T_70_2; // @[Mux.scala 80:57]
  wire [21:0] _T_74_2 = _T_198 ? tagArrayWire_32_2 : _T_72_2; // @[Mux.scala 80:57]
  wire [21:0] _T_76_2 = _T_200 ? tagArrayWire_33_2 : _T_74_2; // @[Mux.scala 80:57]
  wire [21:0] _T_78_2 = _T_202 ? tagArrayWire_34_2 : _T_76_2; // @[Mux.scala 80:57]
  wire [21:0] _T_80_2 = _T_204 ? tagArrayWire_35_2 : _T_78_2; // @[Mux.scala 80:57]
  wire [21:0] _T_82_2 = _T_206 ? tagArrayWire_36_2 : _T_80_2; // @[Mux.scala 80:57]
  wire [21:0] _T_84_2 = _T_208 ? tagArrayWire_37_2 : _T_82_2; // @[Mux.scala 80:57]
  wire [21:0] _T_86_2 = _T_210 ? tagArrayWire_38_2 : _T_84_2; // @[Mux.scala 80:57]
  wire [21:0] _T_88_2 = _T_212 ? tagArrayWire_39_2 : _T_86_2; // @[Mux.scala 80:57]
  wire [21:0] _T_90_2 = _T_214 ? tagArrayWire_40_2 : _T_88_2; // @[Mux.scala 80:57]
  wire [21:0] _T_92_2 = _T_216 ? tagArrayWire_41_2 : _T_90_2; // @[Mux.scala 80:57]
  wire [21:0] _T_94_2 = _T_218 ? tagArrayWire_42_2 : _T_92_2; // @[Mux.scala 80:57]
  wire [21:0] _T_96_2 = _T_220 ? tagArrayWire_43_2 : _T_94_2; // @[Mux.scala 80:57]
  wire [21:0] _T_98_2 = _T_222 ? tagArrayWire_44_2 : _T_96_2; // @[Mux.scala 80:57]
  wire [21:0] _T_100_2 = _T_224 ? tagArrayWire_45_2 : _T_98_2; // @[Mux.scala 80:57]
  wire [21:0] _T_102_2 = _T_226 ? tagArrayWire_46_2 : _T_100_2; // @[Mux.scala 80:57]
  wire [21:0] _T_104_2 = _T_228 ? tagArrayWire_47_2 : _T_102_2; // @[Mux.scala 80:57]
  wire [21:0] _T_106_2 = _T_230 ? tagArrayWire_48_2 : _T_104_2; // @[Mux.scala 80:57]
  wire [21:0] _T_108_2 = _T_232 ? tagArrayWire_49_2 : _T_106_2; // @[Mux.scala 80:57]
  wire [21:0] _T_110_2 = _T_234 ? tagArrayWire_50_2 : _T_108_2; // @[Mux.scala 80:57]
  wire [21:0] _T_112_2 = _T_236 ? tagArrayWire_51_2 : _T_110_2; // @[Mux.scala 80:57]
  wire [21:0] _T_114_2 = _T_238 ? tagArrayWire_52_2 : _T_112_2; // @[Mux.scala 80:57]
  wire [21:0] _T_116_2 = _T_240 ? tagArrayWire_53_2 : _T_114_2; // @[Mux.scala 80:57]
  wire [21:0] _T_118_2 = _T_242 ? tagArrayWire_54_2 : _T_116_2; // @[Mux.scala 80:57]
  wire [21:0] _T_120_2 = _T_244 ? tagArrayWire_55_2 : _T_118_2; // @[Mux.scala 80:57]
  wire [21:0] _T_122_2 = _T_246 ? tagArrayWire_56_2 : _T_120_2; // @[Mux.scala 80:57]
  wire [21:0] _T_124_2 = _T_248 ? tagArrayWire_57_2 : _T_122_2; // @[Mux.scala 80:57]
  wire [21:0] _T_126_2 = _T_250 ? tagArrayWire_58_2 : _T_124_2; // @[Mux.scala 80:57]
  wire [21:0] _T_128_2 = _T_252 ? tagArrayWire_59_2 : _T_126_2; // @[Mux.scala 80:57]
  wire [21:0] _T_130_2 = _T_254 ? tagArrayWire_60_2 : _T_128_2; // @[Mux.scala 80:57]
  wire [21:0] _T_132_2 = _T_256 ? tagArrayWire_61_2 : _T_130_2; // @[Mux.scala 80:57]
  wire [21:0] _T_134_2 = _T_258 ? tagArrayWire_62_2 : _T_132_2; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_2 = _T_260 ? tagArrayWire_63_2 : _T_134_2; // @[Mux.scala 80:57]
  wire  _T_263 = tagMuxOut_2 == tag; // @[Cache.scala 243:76]
  wire  hitArray_2 = vMuxOut_2 & _T_263; // @[Cache.scala 243:60]
  wire  _T_267 = _T_266 | hitArray_2; // @[Cache.scala 244:49]
  reg  vArrayWire_63_3; // @[Reg.scala 27:20]
  reg  vArrayWire_62_3; // @[Reg.scala 27:20]
  reg  vArrayWire_61_3; // @[Reg.scala 27:20]
  reg  vArrayWire_60_3; // @[Reg.scala 27:20]
  reg  vArrayWire_59_3; // @[Reg.scala 27:20]
  reg  vArrayWire_58_3; // @[Reg.scala 27:20]
  reg  vArrayWire_57_3; // @[Reg.scala 27:20]
  reg  vArrayWire_56_3; // @[Reg.scala 27:20]
  reg  vArrayWire_55_3; // @[Reg.scala 27:20]
  reg  vArrayWire_54_3; // @[Reg.scala 27:20]
  reg  vArrayWire_53_3; // @[Reg.scala 27:20]
  reg  vArrayWire_52_3; // @[Reg.scala 27:20]
  reg  vArrayWire_51_3; // @[Reg.scala 27:20]
  reg  vArrayWire_50_3; // @[Reg.scala 27:20]
  reg  vArrayWire_49_3; // @[Reg.scala 27:20]
  reg  vArrayWire_48_3; // @[Reg.scala 27:20]
  reg  vArrayWire_47_3; // @[Reg.scala 27:20]
  reg  vArrayWire_46_3; // @[Reg.scala 27:20]
  reg  vArrayWire_45_3; // @[Reg.scala 27:20]
  reg  vArrayWire_44_3; // @[Reg.scala 27:20]
  reg  vArrayWire_43_3; // @[Reg.scala 27:20]
  reg  vArrayWire_42_3; // @[Reg.scala 27:20]
  reg  vArrayWire_41_3; // @[Reg.scala 27:20]
  reg  vArrayWire_40_3; // @[Reg.scala 27:20]
  reg  vArrayWire_39_3; // @[Reg.scala 27:20]
  reg  vArrayWire_38_3; // @[Reg.scala 27:20]
  reg  vArrayWire_37_3; // @[Reg.scala 27:20]
  reg  vArrayWire_36_3; // @[Reg.scala 27:20]
  reg  vArrayWire_35_3; // @[Reg.scala 27:20]
  reg  vArrayWire_34_3; // @[Reg.scala 27:20]
  reg  vArrayWire_33_3; // @[Reg.scala 27:20]
  reg  vArrayWire_32_3; // @[Reg.scala 27:20]
  reg  vArrayWire_31_3; // @[Reg.scala 27:20]
  reg  vArrayWire_30_3; // @[Reg.scala 27:20]
  reg  vArrayWire_29_3; // @[Reg.scala 27:20]
  reg  vArrayWire_28_3; // @[Reg.scala 27:20]
  reg  vArrayWire_27_3; // @[Reg.scala 27:20]
  reg  vArrayWire_26_3; // @[Reg.scala 27:20]
  reg  vArrayWire_25_3; // @[Reg.scala 27:20]
  reg  vArrayWire_24_3; // @[Reg.scala 27:20]
  reg  vArrayWire_23_3; // @[Reg.scala 27:20]
  reg  vArrayWire_22_3; // @[Reg.scala 27:20]
  reg  vArrayWire_21_3; // @[Reg.scala 27:20]
  reg  vArrayWire_20_3; // @[Reg.scala 27:20]
  reg  vArrayWire_19_3; // @[Reg.scala 27:20]
  reg  vArrayWire_18_3; // @[Reg.scala 27:20]
  reg  vArrayWire_17_3; // @[Reg.scala 27:20]
  reg  vArrayWire_16_3; // @[Reg.scala 27:20]
  reg  vArrayWire_15_3; // @[Reg.scala 27:20]
  reg  vArrayWire_14_3; // @[Reg.scala 27:20]
  reg  vArrayWire_13_3; // @[Reg.scala 27:20]
  reg  vArrayWire_12_3; // @[Reg.scala 27:20]
  reg  vArrayWire_11_3; // @[Reg.scala 27:20]
  reg  vArrayWire_10_3; // @[Reg.scala 27:20]
  reg  vArrayWire_9_3; // @[Reg.scala 27:20]
  reg  vArrayWire_8_3; // @[Reg.scala 27:20]
  reg  vArrayWire_7_3; // @[Reg.scala 27:20]
  reg  vArrayWire_6_3; // @[Reg.scala 27:20]
  reg  vArrayWire_5_3; // @[Reg.scala 27:20]
  reg  vArrayWire_4_3; // @[Reg.scala 27:20]
  reg  vArrayWire_3_3; // @[Reg.scala 27:20]
  reg  vArrayWire_2_3; // @[Reg.scala 27:20]
  reg  vArrayWire_1_3; // @[Reg.scala 27:20]
  reg  vArrayWire_0_3; // @[Reg.scala 27:20]
  wire  _T_137_3 = _T_136 ? vArrayWire_1_3 : vArrayWire_0_3; // @[Mux.scala 80:57]
  wire  _T_139_3 = _T_138 ? vArrayWire_2_3 : _T_137_3; // @[Mux.scala 80:57]
  wire  _T_141_3 = _T_140 ? vArrayWire_3_3 : _T_139_3; // @[Mux.scala 80:57]
  wire  _T_143_3 = _T_142 ? vArrayWire_4_3 : _T_141_3; // @[Mux.scala 80:57]
  wire  _T_145_3 = _T_144 ? vArrayWire_5_3 : _T_143_3; // @[Mux.scala 80:57]
  wire  _T_147_3 = _T_146 ? vArrayWire_6_3 : _T_145_3; // @[Mux.scala 80:57]
  wire  _T_149_3 = _T_148 ? vArrayWire_7_3 : _T_147_3; // @[Mux.scala 80:57]
  wire  _T_151_3 = _T_150 ? vArrayWire_8_3 : _T_149_3; // @[Mux.scala 80:57]
  wire  _T_153_3 = _T_152 ? vArrayWire_9_3 : _T_151_3; // @[Mux.scala 80:57]
  wire  _T_155_3 = _T_154 ? vArrayWire_10_3 : _T_153_3; // @[Mux.scala 80:57]
  wire  _T_157_3 = _T_156 ? vArrayWire_11_3 : _T_155_3; // @[Mux.scala 80:57]
  wire  _T_159_3 = _T_158 ? vArrayWire_12_3 : _T_157_3; // @[Mux.scala 80:57]
  wire  _T_161_3 = _T_160 ? vArrayWire_13_3 : _T_159_3; // @[Mux.scala 80:57]
  wire  _T_163_3 = _T_162 ? vArrayWire_14_3 : _T_161_3; // @[Mux.scala 80:57]
  wire  _T_165_3 = _T_164 ? vArrayWire_15_3 : _T_163_3; // @[Mux.scala 80:57]
  wire  _T_167_3 = _T_166 ? vArrayWire_16_3 : _T_165_3; // @[Mux.scala 80:57]
  wire  _T_169_3 = _T_168 ? vArrayWire_17_3 : _T_167_3; // @[Mux.scala 80:57]
  wire  _T_171_3 = _T_170 ? vArrayWire_18_3 : _T_169_3; // @[Mux.scala 80:57]
  wire  _T_173_3 = _T_172 ? vArrayWire_19_3 : _T_171_3; // @[Mux.scala 80:57]
  wire  _T_175_3 = _T_174 ? vArrayWire_20_3 : _T_173_3; // @[Mux.scala 80:57]
  wire  _T_177_3 = _T_176 ? vArrayWire_21_3 : _T_175_3; // @[Mux.scala 80:57]
  wire  _T_179_3 = _T_178 ? vArrayWire_22_3 : _T_177_3; // @[Mux.scala 80:57]
  wire  _T_181_3 = _T_180 ? vArrayWire_23_3 : _T_179_3; // @[Mux.scala 80:57]
  wire  _T_183_3 = _T_182 ? vArrayWire_24_3 : _T_181_3; // @[Mux.scala 80:57]
  wire  _T_185_3 = _T_184 ? vArrayWire_25_3 : _T_183_3; // @[Mux.scala 80:57]
  wire  _T_187_3 = _T_186 ? vArrayWire_26_3 : _T_185_3; // @[Mux.scala 80:57]
  wire  _T_189_3 = _T_188 ? vArrayWire_27_3 : _T_187_3; // @[Mux.scala 80:57]
  wire  _T_191_3 = _T_190 ? vArrayWire_28_3 : _T_189_3; // @[Mux.scala 80:57]
  wire  _T_193_3 = _T_192 ? vArrayWire_29_3 : _T_191_3; // @[Mux.scala 80:57]
  wire  _T_195_3 = _T_194 ? vArrayWire_30_3 : _T_193_3; // @[Mux.scala 80:57]
  wire  _T_197_3 = _T_196 ? vArrayWire_31_3 : _T_195_3; // @[Mux.scala 80:57]
  wire  _T_199_3 = _T_198 ? vArrayWire_32_3 : _T_197_3; // @[Mux.scala 80:57]
  wire  _T_201_3 = _T_200 ? vArrayWire_33_3 : _T_199_3; // @[Mux.scala 80:57]
  wire  _T_203_3 = _T_202 ? vArrayWire_34_3 : _T_201_3; // @[Mux.scala 80:57]
  wire  _T_205_3 = _T_204 ? vArrayWire_35_3 : _T_203_3; // @[Mux.scala 80:57]
  wire  _T_207_3 = _T_206 ? vArrayWire_36_3 : _T_205_3; // @[Mux.scala 80:57]
  wire  _T_209_3 = _T_208 ? vArrayWire_37_3 : _T_207_3; // @[Mux.scala 80:57]
  wire  _T_211_3 = _T_210 ? vArrayWire_38_3 : _T_209_3; // @[Mux.scala 80:57]
  wire  _T_213_3 = _T_212 ? vArrayWire_39_3 : _T_211_3; // @[Mux.scala 80:57]
  wire  _T_215_3 = _T_214 ? vArrayWire_40_3 : _T_213_3; // @[Mux.scala 80:57]
  wire  _T_217_3 = _T_216 ? vArrayWire_41_3 : _T_215_3; // @[Mux.scala 80:57]
  wire  _T_219_3 = _T_218 ? vArrayWire_42_3 : _T_217_3; // @[Mux.scala 80:57]
  wire  _T_221_3 = _T_220 ? vArrayWire_43_3 : _T_219_3; // @[Mux.scala 80:57]
  wire  _T_223_3 = _T_222 ? vArrayWire_44_3 : _T_221_3; // @[Mux.scala 80:57]
  wire  _T_225_3 = _T_224 ? vArrayWire_45_3 : _T_223_3; // @[Mux.scala 80:57]
  wire  _T_227_3 = _T_226 ? vArrayWire_46_3 : _T_225_3; // @[Mux.scala 80:57]
  wire  _T_229_3 = _T_228 ? vArrayWire_47_3 : _T_227_3; // @[Mux.scala 80:57]
  wire  _T_231_3 = _T_230 ? vArrayWire_48_3 : _T_229_3; // @[Mux.scala 80:57]
  wire  _T_233_3 = _T_232 ? vArrayWire_49_3 : _T_231_3; // @[Mux.scala 80:57]
  wire  _T_235_3 = _T_234 ? vArrayWire_50_3 : _T_233_3; // @[Mux.scala 80:57]
  wire  _T_237_3 = _T_236 ? vArrayWire_51_3 : _T_235_3; // @[Mux.scala 80:57]
  wire  _T_239_3 = _T_238 ? vArrayWire_52_3 : _T_237_3; // @[Mux.scala 80:57]
  wire  _T_241_3 = _T_240 ? vArrayWire_53_3 : _T_239_3; // @[Mux.scala 80:57]
  wire  _T_243_3 = _T_242 ? vArrayWire_54_3 : _T_241_3; // @[Mux.scala 80:57]
  wire  _T_245_3 = _T_244 ? vArrayWire_55_3 : _T_243_3; // @[Mux.scala 80:57]
  wire  _T_247_3 = _T_246 ? vArrayWire_56_3 : _T_245_3; // @[Mux.scala 80:57]
  wire  _T_249_3 = _T_248 ? vArrayWire_57_3 : _T_247_3; // @[Mux.scala 80:57]
  wire  _T_251_3 = _T_250 ? vArrayWire_58_3 : _T_249_3; // @[Mux.scala 80:57]
  wire  _T_253_3 = _T_252 ? vArrayWire_59_3 : _T_251_3; // @[Mux.scala 80:57]
  wire  _T_255_3 = _T_254 ? vArrayWire_60_3 : _T_253_3; // @[Mux.scala 80:57]
  wire  _T_257_3 = _T_256 ? vArrayWire_61_3 : _T_255_3; // @[Mux.scala 80:57]
  wire  _T_259_3 = _T_258 ? vArrayWire_62_3 : _T_257_3; // @[Mux.scala 80:57]
  wire  vMuxOut_3 = _T_260 ? vArrayWire_63_3 : _T_259_3; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_3; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_3; // @[Reg.scala 27:20]
  wire [21:0] _T_12_3 = _T_136 ? tagArrayWire_1_3 : tagArrayWire_0_3; // @[Mux.scala 80:57]
  wire [21:0] _T_14_3 = _T_138 ? tagArrayWire_2_3 : _T_12_3; // @[Mux.scala 80:57]
  wire [21:0] _T_16_3 = _T_140 ? tagArrayWire_3_3 : _T_14_3; // @[Mux.scala 80:57]
  wire [21:0] _T_18_3 = _T_142 ? tagArrayWire_4_3 : _T_16_3; // @[Mux.scala 80:57]
  wire [21:0] _T_20_3 = _T_144 ? tagArrayWire_5_3 : _T_18_3; // @[Mux.scala 80:57]
  wire [21:0] _T_22_3 = _T_146 ? tagArrayWire_6_3 : _T_20_3; // @[Mux.scala 80:57]
  wire [21:0] _T_24_3 = _T_148 ? tagArrayWire_7_3 : _T_22_3; // @[Mux.scala 80:57]
  wire [21:0] _T_26_3 = _T_150 ? tagArrayWire_8_3 : _T_24_3; // @[Mux.scala 80:57]
  wire [21:0] _T_28_3 = _T_152 ? tagArrayWire_9_3 : _T_26_3; // @[Mux.scala 80:57]
  wire [21:0] _T_30_3 = _T_154 ? tagArrayWire_10_3 : _T_28_3; // @[Mux.scala 80:57]
  wire [21:0] _T_32_3 = _T_156 ? tagArrayWire_11_3 : _T_30_3; // @[Mux.scala 80:57]
  wire [21:0] _T_34_3 = _T_158 ? tagArrayWire_12_3 : _T_32_3; // @[Mux.scala 80:57]
  wire [21:0] _T_36_3 = _T_160 ? tagArrayWire_13_3 : _T_34_3; // @[Mux.scala 80:57]
  wire [21:0] _T_38_3 = _T_162 ? tagArrayWire_14_3 : _T_36_3; // @[Mux.scala 80:57]
  wire [21:0] _T_40_3 = _T_164 ? tagArrayWire_15_3 : _T_38_3; // @[Mux.scala 80:57]
  wire [21:0] _T_42_3 = _T_166 ? tagArrayWire_16_3 : _T_40_3; // @[Mux.scala 80:57]
  wire [21:0] _T_44_3 = _T_168 ? tagArrayWire_17_3 : _T_42_3; // @[Mux.scala 80:57]
  wire [21:0] _T_46_3 = _T_170 ? tagArrayWire_18_3 : _T_44_3; // @[Mux.scala 80:57]
  wire [21:0] _T_48_3 = _T_172 ? tagArrayWire_19_3 : _T_46_3; // @[Mux.scala 80:57]
  wire [21:0] _T_50_3 = _T_174 ? tagArrayWire_20_3 : _T_48_3; // @[Mux.scala 80:57]
  wire [21:0] _T_52_3 = _T_176 ? tagArrayWire_21_3 : _T_50_3; // @[Mux.scala 80:57]
  wire [21:0] _T_54_3 = _T_178 ? tagArrayWire_22_3 : _T_52_3; // @[Mux.scala 80:57]
  wire [21:0] _T_56_3 = _T_180 ? tagArrayWire_23_3 : _T_54_3; // @[Mux.scala 80:57]
  wire [21:0] _T_58_3 = _T_182 ? tagArrayWire_24_3 : _T_56_3; // @[Mux.scala 80:57]
  wire [21:0] _T_60_3 = _T_184 ? tagArrayWire_25_3 : _T_58_3; // @[Mux.scala 80:57]
  wire [21:0] _T_62_3 = _T_186 ? tagArrayWire_26_3 : _T_60_3; // @[Mux.scala 80:57]
  wire [21:0] _T_64_3 = _T_188 ? tagArrayWire_27_3 : _T_62_3; // @[Mux.scala 80:57]
  wire [21:0] _T_66_3 = _T_190 ? tagArrayWire_28_3 : _T_64_3; // @[Mux.scala 80:57]
  wire [21:0] _T_68_3 = _T_192 ? tagArrayWire_29_3 : _T_66_3; // @[Mux.scala 80:57]
  wire [21:0] _T_70_3 = _T_194 ? tagArrayWire_30_3 : _T_68_3; // @[Mux.scala 80:57]
  wire [21:0] _T_72_3 = _T_196 ? tagArrayWire_31_3 : _T_70_3; // @[Mux.scala 80:57]
  wire [21:0] _T_74_3 = _T_198 ? tagArrayWire_32_3 : _T_72_3; // @[Mux.scala 80:57]
  wire [21:0] _T_76_3 = _T_200 ? tagArrayWire_33_3 : _T_74_3; // @[Mux.scala 80:57]
  wire [21:0] _T_78_3 = _T_202 ? tagArrayWire_34_3 : _T_76_3; // @[Mux.scala 80:57]
  wire [21:0] _T_80_3 = _T_204 ? tagArrayWire_35_3 : _T_78_3; // @[Mux.scala 80:57]
  wire [21:0] _T_82_3 = _T_206 ? tagArrayWire_36_3 : _T_80_3; // @[Mux.scala 80:57]
  wire [21:0] _T_84_3 = _T_208 ? tagArrayWire_37_3 : _T_82_3; // @[Mux.scala 80:57]
  wire [21:0] _T_86_3 = _T_210 ? tagArrayWire_38_3 : _T_84_3; // @[Mux.scala 80:57]
  wire [21:0] _T_88_3 = _T_212 ? tagArrayWire_39_3 : _T_86_3; // @[Mux.scala 80:57]
  wire [21:0] _T_90_3 = _T_214 ? tagArrayWire_40_3 : _T_88_3; // @[Mux.scala 80:57]
  wire [21:0] _T_92_3 = _T_216 ? tagArrayWire_41_3 : _T_90_3; // @[Mux.scala 80:57]
  wire [21:0] _T_94_3 = _T_218 ? tagArrayWire_42_3 : _T_92_3; // @[Mux.scala 80:57]
  wire [21:0] _T_96_3 = _T_220 ? tagArrayWire_43_3 : _T_94_3; // @[Mux.scala 80:57]
  wire [21:0] _T_98_3 = _T_222 ? tagArrayWire_44_3 : _T_96_3; // @[Mux.scala 80:57]
  wire [21:0] _T_100_3 = _T_224 ? tagArrayWire_45_3 : _T_98_3; // @[Mux.scala 80:57]
  wire [21:0] _T_102_3 = _T_226 ? tagArrayWire_46_3 : _T_100_3; // @[Mux.scala 80:57]
  wire [21:0] _T_104_3 = _T_228 ? tagArrayWire_47_3 : _T_102_3; // @[Mux.scala 80:57]
  wire [21:0] _T_106_3 = _T_230 ? tagArrayWire_48_3 : _T_104_3; // @[Mux.scala 80:57]
  wire [21:0] _T_108_3 = _T_232 ? tagArrayWire_49_3 : _T_106_3; // @[Mux.scala 80:57]
  wire [21:0] _T_110_3 = _T_234 ? tagArrayWire_50_3 : _T_108_3; // @[Mux.scala 80:57]
  wire [21:0] _T_112_3 = _T_236 ? tagArrayWire_51_3 : _T_110_3; // @[Mux.scala 80:57]
  wire [21:0] _T_114_3 = _T_238 ? tagArrayWire_52_3 : _T_112_3; // @[Mux.scala 80:57]
  wire [21:0] _T_116_3 = _T_240 ? tagArrayWire_53_3 : _T_114_3; // @[Mux.scala 80:57]
  wire [21:0] _T_118_3 = _T_242 ? tagArrayWire_54_3 : _T_116_3; // @[Mux.scala 80:57]
  wire [21:0] _T_120_3 = _T_244 ? tagArrayWire_55_3 : _T_118_3; // @[Mux.scala 80:57]
  wire [21:0] _T_122_3 = _T_246 ? tagArrayWire_56_3 : _T_120_3; // @[Mux.scala 80:57]
  wire [21:0] _T_124_3 = _T_248 ? tagArrayWire_57_3 : _T_122_3; // @[Mux.scala 80:57]
  wire [21:0] _T_126_3 = _T_250 ? tagArrayWire_58_3 : _T_124_3; // @[Mux.scala 80:57]
  wire [21:0] _T_128_3 = _T_252 ? tagArrayWire_59_3 : _T_126_3; // @[Mux.scala 80:57]
  wire [21:0] _T_130_3 = _T_254 ? tagArrayWire_60_3 : _T_128_3; // @[Mux.scala 80:57]
  wire [21:0] _T_132_3 = _T_256 ? tagArrayWire_61_3 : _T_130_3; // @[Mux.scala 80:57]
  wire [21:0] _T_134_3 = _T_258 ? tagArrayWire_62_3 : _T_132_3; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_3 = _T_260 ? tagArrayWire_63_3 : _T_134_3; // @[Mux.scala 80:57]
  wire  _T_264 = tagMuxOut_3 == tag; // @[Cache.scala 243:76]
  wire  hitArray_3 = vMuxOut_3 & _T_264; // @[Cache.scala 243:60]
  wire  hit = _T_267 | hitArray_3; // @[Cache.scala 244:49]
  wire  _T_5 = 2'h1 == cacheState; // @[Mux.scala 80:60]
  wire  _T_7 = 2'h2 == cacheState; // @[Mux.scala 80:60]
  wire  _T_9 = 2'h3 == cacheState; // @[Mux.scala 80:60]
  wire  isIdle = cacheState == 2'h0; // @[Cache.scala 214:27]
  wire  isMiss = cacheState == 2'h1; // @[Cache.scala 215:27]
  wire  isWrite = cacheState == 2'h2; // @[Cache.scala 216:28]
  wire  isBlock = cacheState == 2'h3; // @[Cache.scala 217:28]
  wire [127:0] _T_269 = hitArray_0 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_270 = hitArray_1 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_271 = hitArray_2 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_272 = hitArray_3 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _T_273 = _T_269 | _T_270; // @[Mux.scala 27:72]
  wire [127:0] _T_274 = _T_273 | _T_271; // @[Mux.scala 27:72]
  wire [127:0] waysel = _T_274 | _T_272; // @[Mux.scala 27:72]
  reg [1:0] selArrayWire_1; // @[Reg.scala 27:20]
  reg [1:0] selArrayWire_0; // @[Reg.scala 27:20]
  wire [1:0] _T_281 = _T_136 ? selArrayWire_1 : selArrayWire_0; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_2; // @[Reg.scala 27:20]
  wire [1:0] _T_283 = _T_138 ? selArrayWire_2 : _T_281; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_3; // @[Reg.scala 27:20]
  wire [1:0] _T_285 = _T_140 ? selArrayWire_3 : _T_283; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_4; // @[Reg.scala 27:20]
  wire [1:0] _T_287 = _T_142 ? selArrayWire_4 : _T_285; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_5; // @[Reg.scala 27:20]
  wire [1:0] _T_289 = _T_144 ? selArrayWire_5 : _T_287; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_6; // @[Reg.scala 27:20]
  wire [1:0] _T_291 = _T_146 ? selArrayWire_6 : _T_289; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_7; // @[Reg.scala 27:20]
  wire [1:0] _T_293 = _T_148 ? selArrayWire_7 : _T_291; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_8; // @[Reg.scala 27:20]
  wire [1:0] _T_295 = _T_150 ? selArrayWire_8 : _T_293; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_9; // @[Reg.scala 27:20]
  wire [1:0] _T_297 = _T_152 ? selArrayWire_9 : _T_295; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_10; // @[Reg.scala 27:20]
  wire [1:0] _T_299 = _T_154 ? selArrayWire_10 : _T_297; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_11; // @[Reg.scala 27:20]
  wire [1:0] _T_301 = _T_156 ? selArrayWire_11 : _T_299; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_12; // @[Reg.scala 27:20]
  wire [1:0] _T_303 = _T_158 ? selArrayWire_12 : _T_301; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_13; // @[Reg.scala 27:20]
  wire [1:0] _T_305 = _T_160 ? selArrayWire_13 : _T_303; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_14; // @[Reg.scala 27:20]
  wire [1:0] _T_307 = _T_162 ? selArrayWire_14 : _T_305; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_15; // @[Reg.scala 27:20]
  wire [1:0] _T_309 = _T_164 ? selArrayWire_15 : _T_307; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_16; // @[Reg.scala 27:20]
  wire [1:0] _T_311 = _T_166 ? selArrayWire_16 : _T_309; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_17; // @[Reg.scala 27:20]
  wire [1:0] _T_313 = _T_168 ? selArrayWire_17 : _T_311; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_18; // @[Reg.scala 27:20]
  wire [1:0] _T_315 = _T_170 ? selArrayWire_18 : _T_313; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_19; // @[Reg.scala 27:20]
  wire [1:0] _T_317 = _T_172 ? selArrayWire_19 : _T_315; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_20; // @[Reg.scala 27:20]
  wire [1:0] _T_319 = _T_174 ? selArrayWire_20 : _T_317; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_21; // @[Reg.scala 27:20]
  wire [1:0] _T_321 = _T_176 ? selArrayWire_21 : _T_319; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_22; // @[Reg.scala 27:20]
  wire [1:0] _T_323 = _T_178 ? selArrayWire_22 : _T_321; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_23; // @[Reg.scala 27:20]
  wire [1:0] _T_325 = _T_180 ? selArrayWire_23 : _T_323; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_24; // @[Reg.scala 27:20]
  wire [1:0] _T_327 = _T_182 ? selArrayWire_24 : _T_325; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_25; // @[Reg.scala 27:20]
  wire [1:0] _T_329 = _T_184 ? selArrayWire_25 : _T_327; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_26; // @[Reg.scala 27:20]
  wire [1:0] _T_331 = _T_186 ? selArrayWire_26 : _T_329; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_27; // @[Reg.scala 27:20]
  wire [1:0] _T_333 = _T_188 ? selArrayWire_27 : _T_331; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_28; // @[Reg.scala 27:20]
  wire [1:0] _T_335 = _T_190 ? selArrayWire_28 : _T_333; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_29; // @[Reg.scala 27:20]
  wire [1:0] _T_337 = _T_192 ? selArrayWire_29 : _T_335; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_30; // @[Reg.scala 27:20]
  wire [1:0] _T_339 = _T_194 ? selArrayWire_30 : _T_337; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_31; // @[Reg.scala 27:20]
  wire [1:0] _T_341 = _T_196 ? selArrayWire_31 : _T_339; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_32; // @[Reg.scala 27:20]
  wire [1:0] _T_343 = _T_198 ? selArrayWire_32 : _T_341; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_33; // @[Reg.scala 27:20]
  wire [1:0] _T_345 = _T_200 ? selArrayWire_33 : _T_343; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_34; // @[Reg.scala 27:20]
  wire [1:0] _T_347 = _T_202 ? selArrayWire_34 : _T_345; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_35; // @[Reg.scala 27:20]
  wire [1:0] _T_349 = _T_204 ? selArrayWire_35 : _T_347; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_36; // @[Reg.scala 27:20]
  wire [1:0] _T_351 = _T_206 ? selArrayWire_36 : _T_349; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_37; // @[Reg.scala 27:20]
  wire [1:0] _T_353 = _T_208 ? selArrayWire_37 : _T_351; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_38; // @[Reg.scala 27:20]
  wire [1:0] _T_355 = _T_210 ? selArrayWire_38 : _T_353; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_39; // @[Reg.scala 27:20]
  wire [1:0] _T_357 = _T_212 ? selArrayWire_39 : _T_355; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_40; // @[Reg.scala 27:20]
  wire [1:0] _T_359 = _T_214 ? selArrayWire_40 : _T_357; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_41; // @[Reg.scala 27:20]
  wire [1:0] _T_361 = _T_216 ? selArrayWire_41 : _T_359; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_42; // @[Reg.scala 27:20]
  wire [1:0] _T_363 = _T_218 ? selArrayWire_42 : _T_361; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_43; // @[Reg.scala 27:20]
  wire [1:0] _T_365 = _T_220 ? selArrayWire_43 : _T_363; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_44; // @[Reg.scala 27:20]
  wire [1:0] _T_367 = _T_222 ? selArrayWire_44 : _T_365; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_45; // @[Reg.scala 27:20]
  wire [1:0] _T_369 = _T_224 ? selArrayWire_45 : _T_367; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_46; // @[Reg.scala 27:20]
  wire [1:0] _T_371 = _T_226 ? selArrayWire_46 : _T_369; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_47; // @[Reg.scala 27:20]
  wire [1:0] _T_373 = _T_228 ? selArrayWire_47 : _T_371; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_48; // @[Reg.scala 27:20]
  wire [1:0] _T_375 = _T_230 ? selArrayWire_48 : _T_373; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_49; // @[Reg.scala 27:20]
  wire [1:0] _T_377 = _T_232 ? selArrayWire_49 : _T_375; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_50; // @[Reg.scala 27:20]
  wire [1:0] _T_379 = _T_234 ? selArrayWire_50 : _T_377; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_51; // @[Reg.scala 27:20]
  wire [1:0] _T_381 = _T_236 ? selArrayWire_51 : _T_379; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_52; // @[Reg.scala 27:20]
  wire [1:0] _T_383 = _T_238 ? selArrayWire_52 : _T_381; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_53; // @[Reg.scala 27:20]
  wire [1:0] _T_385 = _T_240 ? selArrayWire_53 : _T_383; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_54; // @[Reg.scala 27:20]
  wire [1:0] _T_387 = _T_242 ? selArrayWire_54 : _T_385; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_55; // @[Reg.scala 27:20]
  wire [1:0] _T_389 = _T_244 ? selArrayWire_55 : _T_387; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_56; // @[Reg.scala 27:20]
  wire [1:0] _T_391 = _T_246 ? selArrayWire_56 : _T_389; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_57; // @[Reg.scala 27:20]
  wire [1:0] _T_393 = _T_248 ? selArrayWire_57 : _T_391; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_58; // @[Reg.scala 27:20]
  wire [1:0] _T_395 = _T_250 ? selArrayWire_58 : _T_393; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_59; // @[Reg.scala 27:20]
  wire [1:0] _T_397 = _T_252 ? selArrayWire_59 : _T_395; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_60; // @[Reg.scala 27:20]
  wire [1:0] _T_399 = _T_254 ? selArrayWire_60 : _T_397; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_61; // @[Reg.scala 27:20]
  wire [1:0] _T_401 = _T_256 ? selArrayWire_61 : _T_399; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_62; // @[Reg.scala 27:20]
  wire [1:0] _T_403 = _T_258 ? selArrayWire_62 : _T_401; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_63; // @[Reg.scala 27:20]
  wire [1:0] sramSel = _T_260 ? selArrayWire_63 : _T_403; // @[Mux.scala 80:57]
  wire [1:0] _T_408 = selArrayWire_0 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_409 = 6'h0 == index; // @[Cache.scala 292:36]
  wire  _T_410 = io_cacheOut_r_last_i & _T_409; // @[Cache.scala 292:28]
  wire  _T_414 = selArrayWire_0 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_415 = _T_410 & _T_414; // @[Cache.scala 295:85]
  wire  _T_416 = _T_415 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_2 = _T_416 | vArrayWire_0_0; // @[Reg.scala 28:19]
  wire  _T_426 = selArrayWire_0 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_427 = _T_410 & _T_426; // @[Cache.scala 295:85]
  wire  _T_428 = _T_427 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_4 = _T_428 | vArrayWire_0_1; // @[Reg.scala 28:19]
  wire  _T_438 = selArrayWire_0 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_439 = _T_410 & _T_438; // @[Cache.scala 295:85]
  wire  _T_440 = _T_439 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_6 = _T_440 | vArrayWire_0_2; // @[Reg.scala 28:19]
  wire  _T_450 = selArrayWire_0 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_451 = _T_410 & _T_450; // @[Cache.scala 295:85]
  wire  _T_452 = _T_451 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_8 = _T_452 | vArrayWire_0_3; // @[Reg.scala 28:19]
  wire [1:0] _T_461 = selArrayWire_1 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_463 = io_cacheOut_r_last_i & _T_136; // @[Cache.scala 292:28]
  wire  _T_467 = selArrayWire_1 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_468 = _T_463 & _T_467; // @[Cache.scala 295:85]
  wire  _T_469 = _T_468 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_11 = _T_469 | vArrayWire_1_0; // @[Reg.scala 28:19]
  wire  _T_479 = selArrayWire_1 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_480 = _T_463 & _T_479; // @[Cache.scala 295:85]
  wire  _T_481 = _T_480 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_13 = _T_481 | vArrayWire_1_1; // @[Reg.scala 28:19]
  wire  _T_491 = selArrayWire_1 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_492 = _T_463 & _T_491; // @[Cache.scala 295:85]
  wire  _T_493 = _T_492 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_15 = _T_493 | vArrayWire_1_2; // @[Reg.scala 28:19]
  wire  _T_503 = selArrayWire_1 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_504 = _T_463 & _T_503; // @[Cache.scala 295:85]
  wire  _T_505 = _T_504 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_17 = _T_505 | vArrayWire_1_3; // @[Reg.scala 28:19]
  wire [1:0] _T_514 = selArrayWire_2 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_516 = io_cacheOut_r_last_i & _T_138; // @[Cache.scala 292:28]
  wire  _T_520 = selArrayWire_2 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_521 = _T_516 & _T_520; // @[Cache.scala 295:85]
  wire  _T_522 = _T_521 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_20 = _T_522 | vArrayWire_2_0; // @[Reg.scala 28:19]
  wire  _T_532 = selArrayWire_2 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_533 = _T_516 & _T_532; // @[Cache.scala 295:85]
  wire  _T_534 = _T_533 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_22 = _T_534 | vArrayWire_2_1; // @[Reg.scala 28:19]
  wire  _T_544 = selArrayWire_2 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_545 = _T_516 & _T_544; // @[Cache.scala 295:85]
  wire  _T_546 = _T_545 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_24 = _T_546 | vArrayWire_2_2; // @[Reg.scala 28:19]
  wire  _T_556 = selArrayWire_2 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_557 = _T_516 & _T_556; // @[Cache.scala 295:85]
  wire  _T_558 = _T_557 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_26 = _T_558 | vArrayWire_2_3; // @[Reg.scala 28:19]
  wire [1:0] _T_567 = selArrayWire_3 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_569 = io_cacheOut_r_last_i & _T_140; // @[Cache.scala 292:28]
  wire  _T_573 = selArrayWire_3 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_574 = _T_569 & _T_573; // @[Cache.scala 295:85]
  wire  _T_575 = _T_574 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_29 = _T_575 | vArrayWire_3_0; // @[Reg.scala 28:19]
  wire  _T_585 = selArrayWire_3 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_586 = _T_569 & _T_585; // @[Cache.scala 295:85]
  wire  _T_587 = _T_586 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_31 = _T_587 | vArrayWire_3_1; // @[Reg.scala 28:19]
  wire  _T_597 = selArrayWire_3 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_598 = _T_569 & _T_597; // @[Cache.scala 295:85]
  wire  _T_599 = _T_598 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_33 = _T_599 | vArrayWire_3_2; // @[Reg.scala 28:19]
  wire  _T_609 = selArrayWire_3 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_610 = _T_569 & _T_609; // @[Cache.scala 295:85]
  wire  _T_611 = _T_610 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_35 = _T_611 | vArrayWire_3_3; // @[Reg.scala 28:19]
  wire [1:0] _T_620 = selArrayWire_4 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_622 = io_cacheOut_r_last_i & _T_142; // @[Cache.scala 292:28]
  wire  _T_626 = selArrayWire_4 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_627 = _T_622 & _T_626; // @[Cache.scala 295:85]
  wire  _T_628 = _T_627 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_38 = _T_628 | vArrayWire_4_0; // @[Reg.scala 28:19]
  wire  _T_638 = selArrayWire_4 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_639 = _T_622 & _T_638; // @[Cache.scala 295:85]
  wire  _T_640 = _T_639 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_40 = _T_640 | vArrayWire_4_1; // @[Reg.scala 28:19]
  wire  _T_650 = selArrayWire_4 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_651 = _T_622 & _T_650; // @[Cache.scala 295:85]
  wire  _T_652 = _T_651 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_42 = _T_652 | vArrayWire_4_2; // @[Reg.scala 28:19]
  wire  _T_662 = selArrayWire_4 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_663 = _T_622 & _T_662; // @[Cache.scala 295:85]
  wire  _T_664 = _T_663 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_44 = _T_664 | vArrayWire_4_3; // @[Reg.scala 28:19]
  wire [1:0] _T_673 = selArrayWire_5 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_675 = io_cacheOut_r_last_i & _T_144; // @[Cache.scala 292:28]
  wire  _T_679 = selArrayWire_5 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_680 = _T_675 & _T_679; // @[Cache.scala 295:85]
  wire  _T_681 = _T_680 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_47 = _T_681 | vArrayWire_5_0; // @[Reg.scala 28:19]
  wire  _T_691 = selArrayWire_5 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_692 = _T_675 & _T_691; // @[Cache.scala 295:85]
  wire  _T_693 = _T_692 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_49 = _T_693 | vArrayWire_5_1; // @[Reg.scala 28:19]
  wire  _T_703 = selArrayWire_5 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_704 = _T_675 & _T_703; // @[Cache.scala 295:85]
  wire  _T_705 = _T_704 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_51 = _T_705 | vArrayWire_5_2; // @[Reg.scala 28:19]
  wire  _T_715 = selArrayWire_5 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_716 = _T_675 & _T_715; // @[Cache.scala 295:85]
  wire  _T_717 = _T_716 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_53 = _T_717 | vArrayWire_5_3; // @[Reg.scala 28:19]
  wire [1:0] _T_726 = selArrayWire_6 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_728 = io_cacheOut_r_last_i & _T_146; // @[Cache.scala 292:28]
  wire  _T_732 = selArrayWire_6 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_733 = _T_728 & _T_732; // @[Cache.scala 295:85]
  wire  _T_734 = _T_733 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_56 = _T_734 | vArrayWire_6_0; // @[Reg.scala 28:19]
  wire  _T_744 = selArrayWire_6 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_745 = _T_728 & _T_744; // @[Cache.scala 295:85]
  wire  _T_746 = _T_745 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_58 = _T_746 | vArrayWire_6_1; // @[Reg.scala 28:19]
  wire  _T_756 = selArrayWire_6 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_757 = _T_728 & _T_756; // @[Cache.scala 295:85]
  wire  _T_758 = _T_757 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_60 = _T_758 | vArrayWire_6_2; // @[Reg.scala 28:19]
  wire  _T_768 = selArrayWire_6 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_769 = _T_728 & _T_768; // @[Cache.scala 295:85]
  wire  _T_770 = _T_769 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_62 = _T_770 | vArrayWire_6_3; // @[Reg.scala 28:19]
  wire [1:0] _T_779 = selArrayWire_7 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_781 = io_cacheOut_r_last_i & _T_148; // @[Cache.scala 292:28]
  wire  _T_785 = selArrayWire_7 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_786 = _T_781 & _T_785; // @[Cache.scala 295:85]
  wire  _T_787 = _T_786 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_65 = _T_787 | vArrayWire_7_0; // @[Reg.scala 28:19]
  wire  _T_797 = selArrayWire_7 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_798 = _T_781 & _T_797; // @[Cache.scala 295:85]
  wire  _T_799 = _T_798 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_67 = _T_799 | vArrayWire_7_1; // @[Reg.scala 28:19]
  wire  _T_809 = selArrayWire_7 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_810 = _T_781 & _T_809; // @[Cache.scala 295:85]
  wire  _T_811 = _T_810 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_69 = _T_811 | vArrayWire_7_2; // @[Reg.scala 28:19]
  wire  _T_821 = selArrayWire_7 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_822 = _T_781 & _T_821; // @[Cache.scala 295:85]
  wire  _T_823 = _T_822 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_71 = _T_823 | vArrayWire_7_3; // @[Reg.scala 28:19]
  wire [1:0] _T_832 = selArrayWire_8 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_834 = io_cacheOut_r_last_i & _T_150; // @[Cache.scala 292:28]
  wire  _T_838 = selArrayWire_8 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_839 = _T_834 & _T_838; // @[Cache.scala 295:85]
  wire  _T_840 = _T_839 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_74 = _T_840 | vArrayWire_8_0; // @[Reg.scala 28:19]
  wire  _T_850 = selArrayWire_8 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_851 = _T_834 & _T_850; // @[Cache.scala 295:85]
  wire  _T_852 = _T_851 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_76 = _T_852 | vArrayWire_8_1; // @[Reg.scala 28:19]
  wire  _T_862 = selArrayWire_8 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_863 = _T_834 & _T_862; // @[Cache.scala 295:85]
  wire  _T_864 = _T_863 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_78 = _T_864 | vArrayWire_8_2; // @[Reg.scala 28:19]
  wire  _T_874 = selArrayWire_8 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_875 = _T_834 & _T_874; // @[Cache.scala 295:85]
  wire  _T_876 = _T_875 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_80 = _T_876 | vArrayWire_8_3; // @[Reg.scala 28:19]
  wire [1:0] _T_885 = selArrayWire_9 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_887 = io_cacheOut_r_last_i & _T_152; // @[Cache.scala 292:28]
  wire  _T_891 = selArrayWire_9 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_892 = _T_887 & _T_891; // @[Cache.scala 295:85]
  wire  _T_893 = _T_892 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_83 = _T_893 | vArrayWire_9_0; // @[Reg.scala 28:19]
  wire  _T_903 = selArrayWire_9 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_904 = _T_887 & _T_903; // @[Cache.scala 295:85]
  wire  _T_905 = _T_904 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_85 = _T_905 | vArrayWire_9_1; // @[Reg.scala 28:19]
  wire  _T_915 = selArrayWire_9 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_916 = _T_887 & _T_915; // @[Cache.scala 295:85]
  wire  _T_917 = _T_916 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_87 = _T_917 | vArrayWire_9_2; // @[Reg.scala 28:19]
  wire  _T_927 = selArrayWire_9 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_928 = _T_887 & _T_927; // @[Cache.scala 295:85]
  wire  _T_929 = _T_928 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_89 = _T_929 | vArrayWire_9_3; // @[Reg.scala 28:19]
  wire [1:0] _T_938 = selArrayWire_10 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_940 = io_cacheOut_r_last_i & _T_154; // @[Cache.scala 292:28]
  wire  _T_944 = selArrayWire_10 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_945 = _T_940 & _T_944; // @[Cache.scala 295:85]
  wire  _T_946 = _T_945 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_92 = _T_946 | vArrayWire_10_0; // @[Reg.scala 28:19]
  wire  _T_956 = selArrayWire_10 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_957 = _T_940 & _T_956; // @[Cache.scala 295:85]
  wire  _T_958 = _T_957 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_94 = _T_958 | vArrayWire_10_1; // @[Reg.scala 28:19]
  wire  _T_968 = selArrayWire_10 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_969 = _T_940 & _T_968; // @[Cache.scala 295:85]
  wire  _T_970 = _T_969 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_96 = _T_970 | vArrayWire_10_2; // @[Reg.scala 28:19]
  wire  _T_980 = selArrayWire_10 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_981 = _T_940 & _T_980; // @[Cache.scala 295:85]
  wire  _T_982 = _T_981 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_98 = _T_982 | vArrayWire_10_3; // @[Reg.scala 28:19]
  wire [1:0] _T_991 = selArrayWire_11 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_993 = io_cacheOut_r_last_i & _T_156; // @[Cache.scala 292:28]
  wire  _T_997 = selArrayWire_11 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_998 = _T_993 & _T_997; // @[Cache.scala 295:85]
  wire  _T_999 = _T_998 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_101 = _T_999 | vArrayWire_11_0; // @[Reg.scala 28:19]
  wire  _T_1009 = selArrayWire_11 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1010 = _T_993 & _T_1009; // @[Cache.scala 295:85]
  wire  _T_1011 = _T_1010 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_103 = _T_1011 | vArrayWire_11_1; // @[Reg.scala 28:19]
  wire  _T_1021 = selArrayWire_11 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1022 = _T_993 & _T_1021; // @[Cache.scala 295:85]
  wire  _T_1023 = _T_1022 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_105 = _T_1023 | vArrayWire_11_2; // @[Reg.scala 28:19]
  wire  _T_1033 = selArrayWire_11 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1034 = _T_993 & _T_1033; // @[Cache.scala 295:85]
  wire  _T_1035 = _T_1034 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_107 = _T_1035 | vArrayWire_11_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1044 = selArrayWire_12 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1046 = io_cacheOut_r_last_i & _T_158; // @[Cache.scala 292:28]
  wire  _T_1050 = selArrayWire_12 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1051 = _T_1046 & _T_1050; // @[Cache.scala 295:85]
  wire  _T_1052 = _T_1051 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_110 = _T_1052 | vArrayWire_12_0; // @[Reg.scala 28:19]
  wire  _T_1062 = selArrayWire_12 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1063 = _T_1046 & _T_1062; // @[Cache.scala 295:85]
  wire  _T_1064 = _T_1063 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_112 = _T_1064 | vArrayWire_12_1; // @[Reg.scala 28:19]
  wire  _T_1074 = selArrayWire_12 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1075 = _T_1046 & _T_1074; // @[Cache.scala 295:85]
  wire  _T_1076 = _T_1075 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_114 = _T_1076 | vArrayWire_12_2; // @[Reg.scala 28:19]
  wire  _T_1086 = selArrayWire_12 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1087 = _T_1046 & _T_1086; // @[Cache.scala 295:85]
  wire  _T_1088 = _T_1087 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_116 = _T_1088 | vArrayWire_12_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1097 = selArrayWire_13 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1099 = io_cacheOut_r_last_i & _T_160; // @[Cache.scala 292:28]
  wire  _T_1103 = selArrayWire_13 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1104 = _T_1099 & _T_1103; // @[Cache.scala 295:85]
  wire  _T_1105 = _T_1104 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_119 = _T_1105 | vArrayWire_13_0; // @[Reg.scala 28:19]
  wire  _T_1115 = selArrayWire_13 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1116 = _T_1099 & _T_1115; // @[Cache.scala 295:85]
  wire  _T_1117 = _T_1116 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_121 = _T_1117 | vArrayWire_13_1; // @[Reg.scala 28:19]
  wire  _T_1127 = selArrayWire_13 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1128 = _T_1099 & _T_1127; // @[Cache.scala 295:85]
  wire  _T_1129 = _T_1128 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_123 = _T_1129 | vArrayWire_13_2; // @[Reg.scala 28:19]
  wire  _T_1139 = selArrayWire_13 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1140 = _T_1099 & _T_1139; // @[Cache.scala 295:85]
  wire  _T_1141 = _T_1140 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_125 = _T_1141 | vArrayWire_13_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1150 = selArrayWire_14 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1152 = io_cacheOut_r_last_i & _T_162; // @[Cache.scala 292:28]
  wire  _T_1156 = selArrayWire_14 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1157 = _T_1152 & _T_1156; // @[Cache.scala 295:85]
  wire  _T_1158 = _T_1157 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_128 = _T_1158 | vArrayWire_14_0; // @[Reg.scala 28:19]
  wire  _T_1168 = selArrayWire_14 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1169 = _T_1152 & _T_1168; // @[Cache.scala 295:85]
  wire  _T_1170 = _T_1169 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_130 = _T_1170 | vArrayWire_14_1; // @[Reg.scala 28:19]
  wire  _T_1180 = selArrayWire_14 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1181 = _T_1152 & _T_1180; // @[Cache.scala 295:85]
  wire  _T_1182 = _T_1181 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_132 = _T_1182 | vArrayWire_14_2; // @[Reg.scala 28:19]
  wire  _T_1192 = selArrayWire_14 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1193 = _T_1152 & _T_1192; // @[Cache.scala 295:85]
  wire  _T_1194 = _T_1193 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_134 = _T_1194 | vArrayWire_14_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1203 = selArrayWire_15 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1205 = io_cacheOut_r_last_i & _T_164; // @[Cache.scala 292:28]
  wire  _T_1209 = selArrayWire_15 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1210 = _T_1205 & _T_1209; // @[Cache.scala 295:85]
  wire  _T_1211 = _T_1210 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_137 = _T_1211 | vArrayWire_15_0; // @[Reg.scala 28:19]
  wire  _T_1221 = selArrayWire_15 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1222 = _T_1205 & _T_1221; // @[Cache.scala 295:85]
  wire  _T_1223 = _T_1222 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_139 = _T_1223 | vArrayWire_15_1; // @[Reg.scala 28:19]
  wire  _T_1233 = selArrayWire_15 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1234 = _T_1205 & _T_1233; // @[Cache.scala 295:85]
  wire  _T_1235 = _T_1234 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_141 = _T_1235 | vArrayWire_15_2; // @[Reg.scala 28:19]
  wire  _T_1245 = selArrayWire_15 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1246 = _T_1205 & _T_1245; // @[Cache.scala 295:85]
  wire  _T_1247 = _T_1246 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_143 = _T_1247 | vArrayWire_15_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1256 = selArrayWire_16 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1258 = io_cacheOut_r_last_i & _T_166; // @[Cache.scala 292:28]
  wire  _T_1262 = selArrayWire_16 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1263 = _T_1258 & _T_1262; // @[Cache.scala 295:85]
  wire  _T_1264 = _T_1263 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_146 = _T_1264 | vArrayWire_16_0; // @[Reg.scala 28:19]
  wire  _T_1274 = selArrayWire_16 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1275 = _T_1258 & _T_1274; // @[Cache.scala 295:85]
  wire  _T_1276 = _T_1275 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_148 = _T_1276 | vArrayWire_16_1; // @[Reg.scala 28:19]
  wire  _T_1286 = selArrayWire_16 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1287 = _T_1258 & _T_1286; // @[Cache.scala 295:85]
  wire  _T_1288 = _T_1287 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_150 = _T_1288 | vArrayWire_16_2; // @[Reg.scala 28:19]
  wire  _T_1298 = selArrayWire_16 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1299 = _T_1258 & _T_1298; // @[Cache.scala 295:85]
  wire  _T_1300 = _T_1299 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_152 = _T_1300 | vArrayWire_16_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1309 = selArrayWire_17 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1311 = io_cacheOut_r_last_i & _T_168; // @[Cache.scala 292:28]
  wire  _T_1315 = selArrayWire_17 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1316 = _T_1311 & _T_1315; // @[Cache.scala 295:85]
  wire  _T_1317 = _T_1316 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_155 = _T_1317 | vArrayWire_17_0; // @[Reg.scala 28:19]
  wire  _T_1327 = selArrayWire_17 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1328 = _T_1311 & _T_1327; // @[Cache.scala 295:85]
  wire  _T_1329 = _T_1328 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_157 = _T_1329 | vArrayWire_17_1; // @[Reg.scala 28:19]
  wire  _T_1339 = selArrayWire_17 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1340 = _T_1311 & _T_1339; // @[Cache.scala 295:85]
  wire  _T_1341 = _T_1340 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_159 = _T_1341 | vArrayWire_17_2; // @[Reg.scala 28:19]
  wire  _T_1351 = selArrayWire_17 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1352 = _T_1311 & _T_1351; // @[Cache.scala 295:85]
  wire  _T_1353 = _T_1352 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_161 = _T_1353 | vArrayWire_17_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1362 = selArrayWire_18 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1364 = io_cacheOut_r_last_i & _T_170; // @[Cache.scala 292:28]
  wire  _T_1368 = selArrayWire_18 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1369 = _T_1364 & _T_1368; // @[Cache.scala 295:85]
  wire  _T_1370 = _T_1369 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_164 = _T_1370 | vArrayWire_18_0; // @[Reg.scala 28:19]
  wire  _T_1380 = selArrayWire_18 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1381 = _T_1364 & _T_1380; // @[Cache.scala 295:85]
  wire  _T_1382 = _T_1381 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_166 = _T_1382 | vArrayWire_18_1; // @[Reg.scala 28:19]
  wire  _T_1392 = selArrayWire_18 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1393 = _T_1364 & _T_1392; // @[Cache.scala 295:85]
  wire  _T_1394 = _T_1393 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_168 = _T_1394 | vArrayWire_18_2; // @[Reg.scala 28:19]
  wire  _T_1404 = selArrayWire_18 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1405 = _T_1364 & _T_1404; // @[Cache.scala 295:85]
  wire  _T_1406 = _T_1405 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_170 = _T_1406 | vArrayWire_18_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1415 = selArrayWire_19 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1417 = io_cacheOut_r_last_i & _T_172; // @[Cache.scala 292:28]
  wire  _T_1421 = selArrayWire_19 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1422 = _T_1417 & _T_1421; // @[Cache.scala 295:85]
  wire  _T_1423 = _T_1422 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_173 = _T_1423 | vArrayWire_19_0; // @[Reg.scala 28:19]
  wire  _T_1433 = selArrayWire_19 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1434 = _T_1417 & _T_1433; // @[Cache.scala 295:85]
  wire  _T_1435 = _T_1434 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_175 = _T_1435 | vArrayWire_19_1; // @[Reg.scala 28:19]
  wire  _T_1445 = selArrayWire_19 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1446 = _T_1417 & _T_1445; // @[Cache.scala 295:85]
  wire  _T_1447 = _T_1446 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_177 = _T_1447 | vArrayWire_19_2; // @[Reg.scala 28:19]
  wire  _T_1457 = selArrayWire_19 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1458 = _T_1417 & _T_1457; // @[Cache.scala 295:85]
  wire  _T_1459 = _T_1458 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_179 = _T_1459 | vArrayWire_19_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1468 = selArrayWire_20 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1470 = io_cacheOut_r_last_i & _T_174; // @[Cache.scala 292:28]
  wire  _T_1474 = selArrayWire_20 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1475 = _T_1470 & _T_1474; // @[Cache.scala 295:85]
  wire  _T_1476 = _T_1475 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_182 = _T_1476 | vArrayWire_20_0; // @[Reg.scala 28:19]
  wire  _T_1486 = selArrayWire_20 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1487 = _T_1470 & _T_1486; // @[Cache.scala 295:85]
  wire  _T_1488 = _T_1487 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_184 = _T_1488 | vArrayWire_20_1; // @[Reg.scala 28:19]
  wire  _T_1498 = selArrayWire_20 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1499 = _T_1470 & _T_1498; // @[Cache.scala 295:85]
  wire  _T_1500 = _T_1499 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_186 = _T_1500 | vArrayWire_20_2; // @[Reg.scala 28:19]
  wire  _T_1510 = selArrayWire_20 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1511 = _T_1470 & _T_1510; // @[Cache.scala 295:85]
  wire  _T_1512 = _T_1511 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_188 = _T_1512 | vArrayWire_20_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1521 = selArrayWire_21 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1523 = io_cacheOut_r_last_i & _T_176; // @[Cache.scala 292:28]
  wire  _T_1527 = selArrayWire_21 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1528 = _T_1523 & _T_1527; // @[Cache.scala 295:85]
  wire  _T_1529 = _T_1528 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_191 = _T_1529 | vArrayWire_21_0; // @[Reg.scala 28:19]
  wire  _T_1539 = selArrayWire_21 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1540 = _T_1523 & _T_1539; // @[Cache.scala 295:85]
  wire  _T_1541 = _T_1540 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_193 = _T_1541 | vArrayWire_21_1; // @[Reg.scala 28:19]
  wire  _T_1551 = selArrayWire_21 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1552 = _T_1523 & _T_1551; // @[Cache.scala 295:85]
  wire  _T_1553 = _T_1552 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_195 = _T_1553 | vArrayWire_21_2; // @[Reg.scala 28:19]
  wire  _T_1563 = selArrayWire_21 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1564 = _T_1523 & _T_1563; // @[Cache.scala 295:85]
  wire  _T_1565 = _T_1564 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_197 = _T_1565 | vArrayWire_21_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1574 = selArrayWire_22 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1576 = io_cacheOut_r_last_i & _T_178; // @[Cache.scala 292:28]
  wire  _T_1580 = selArrayWire_22 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1581 = _T_1576 & _T_1580; // @[Cache.scala 295:85]
  wire  _T_1582 = _T_1581 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_200 = _T_1582 | vArrayWire_22_0; // @[Reg.scala 28:19]
  wire  _T_1592 = selArrayWire_22 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1593 = _T_1576 & _T_1592; // @[Cache.scala 295:85]
  wire  _T_1594 = _T_1593 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_202 = _T_1594 | vArrayWire_22_1; // @[Reg.scala 28:19]
  wire  _T_1604 = selArrayWire_22 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1605 = _T_1576 & _T_1604; // @[Cache.scala 295:85]
  wire  _T_1606 = _T_1605 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_204 = _T_1606 | vArrayWire_22_2; // @[Reg.scala 28:19]
  wire  _T_1616 = selArrayWire_22 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1617 = _T_1576 & _T_1616; // @[Cache.scala 295:85]
  wire  _T_1618 = _T_1617 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_206 = _T_1618 | vArrayWire_22_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1627 = selArrayWire_23 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1629 = io_cacheOut_r_last_i & _T_180; // @[Cache.scala 292:28]
  wire  _T_1633 = selArrayWire_23 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1634 = _T_1629 & _T_1633; // @[Cache.scala 295:85]
  wire  _T_1635 = _T_1634 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_209 = _T_1635 | vArrayWire_23_0; // @[Reg.scala 28:19]
  wire  _T_1645 = selArrayWire_23 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1646 = _T_1629 & _T_1645; // @[Cache.scala 295:85]
  wire  _T_1647 = _T_1646 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_211 = _T_1647 | vArrayWire_23_1; // @[Reg.scala 28:19]
  wire  _T_1657 = selArrayWire_23 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1658 = _T_1629 & _T_1657; // @[Cache.scala 295:85]
  wire  _T_1659 = _T_1658 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_213 = _T_1659 | vArrayWire_23_2; // @[Reg.scala 28:19]
  wire  _T_1669 = selArrayWire_23 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1670 = _T_1629 & _T_1669; // @[Cache.scala 295:85]
  wire  _T_1671 = _T_1670 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_215 = _T_1671 | vArrayWire_23_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1680 = selArrayWire_24 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1682 = io_cacheOut_r_last_i & _T_182; // @[Cache.scala 292:28]
  wire  _T_1686 = selArrayWire_24 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1687 = _T_1682 & _T_1686; // @[Cache.scala 295:85]
  wire  _T_1688 = _T_1687 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_218 = _T_1688 | vArrayWire_24_0; // @[Reg.scala 28:19]
  wire  _T_1698 = selArrayWire_24 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1699 = _T_1682 & _T_1698; // @[Cache.scala 295:85]
  wire  _T_1700 = _T_1699 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_220 = _T_1700 | vArrayWire_24_1; // @[Reg.scala 28:19]
  wire  _T_1710 = selArrayWire_24 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1711 = _T_1682 & _T_1710; // @[Cache.scala 295:85]
  wire  _T_1712 = _T_1711 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_222 = _T_1712 | vArrayWire_24_2; // @[Reg.scala 28:19]
  wire  _T_1722 = selArrayWire_24 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1723 = _T_1682 & _T_1722; // @[Cache.scala 295:85]
  wire  _T_1724 = _T_1723 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_224 = _T_1724 | vArrayWire_24_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1733 = selArrayWire_25 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1735 = io_cacheOut_r_last_i & _T_184; // @[Cache.scala 292:28]
  wire  _T_1739 = selArrayWire_25 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1740 = _T_1735 & _T_1739; // @[Cache.scala 295:85]
  wire  _T_1741 = _T_1740 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_227 = _T_1741 | vArrayWire_25_0; // @[Reg.scala 28:19]
  wire  _T_1751 = selArrayWire_25 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1752 = _T_1735 & _T_1751; // @[Cache.scala 295:85]
  wire  _T_1753 = _T_1752 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_229 = _T_1753 | vArrayWire_25_1; // @[Reg.scala 28:19]
  wire  _T_1763 = selArrayWire_25 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1764 = _T_1735 & _T_1763; // @[Cache.scala 295:85]
  wire  _T_1765 = _T_1764 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_231 = _T_1765 | vArrayWire_25_2; // @[Reg.scala 28:19]
  wire  _T_1775 = selArrayWire_25 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1776 = _T_1735 & _T_1775; // @[Cache.scala 295:85]
  wire  _T_1777 = _T_1776 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_233 = _T_1777 | vArrayWire_25_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1786 = selArrayWire_26 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1788 = io_cacheOut_r_last_i & _T_186; // @[Cache.scala 292:28]
  wire  _T_1792 = selArrayWire_26 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1793 = _T_1788 & _T_1792; // @[Cache.scala 295:85]
  wire  _T_1794 = _T_1793 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_236 = _T_1794 | vArrayWire_26_0; // @[Reg.scala 28:19]
  wire  _T_1804 = selArrayWire_26 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1805 = _T_1788 & _T_1804; // @[Cache.scala 295:85]
  wire  _T_1806 = _T_1805 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_238 = _T_1806 | vArrayWire_26_1; // @[Reg.scala 28:19]
  wire  _T_1816 = selArrayWire_26 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1817 = _T_1788 & _T_1816; // @[Cache.scala 295:85]
  wire  _T_1818 = _T_1817 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_240 = _T_1818 | vArrayWire_26_2; // @[Reg.scala 28:19]
  wire  _T_1828 = selArrayWire_26 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1829 = _T_1788 & _T_1828; // @[Cache.scala 295:85]
  wire  _T_1830 = _T_1829 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_242 = _T_1830 | vArrayWire_26_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1839 = selArrayWire_27 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1841 = io_cacheOut_r_last_i & _T_188; // @[Cache.scala 292:28]
  wire  _T_1845 = selArrayWire_27 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1846 = _T_1841 & _T_1845; // @[Cache.scala 295:85]
  wire  _T_1847 = _T_1846 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_245 = _T_1847 | vArrayWire_27_0; // @[Reg.scala 28:19]
  wire  _T_1857 = selArrayWire_27 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1858 = _T_1841 & _T_1857; // @[Cache.scala 295:85]
  wire  _T_1859 = _T_1858 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_247 = _T_1859 | vArrayWire_27_1; // @[Reg.scala 28:19]
  wire  _T_1869 = selArrayWire_27 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1870 = _T_1841 & _T_1869; // @[Cache.scala 295:85]
  wire  _T_1871 = _T_1870 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_249 = _T_1871 | vArrayWire_27_2; // @[Reg.scala 28:19]
  wire  _T_1881 = selArrayWire_27 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1882 = _T_1841 & _T_1881; // @[Cache.scala 295:85]
  wire  _T_1883 = _T_1882 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_251 = _T_1883 | vArrayWire_27_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1892 = selArrayWire_28 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1894 = io_cacheOut_r_last_i & _T_190; // @[Cache.scala 292:28]
  wire  _T_1898 = selArrayWire_28 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1899 = _T_1894 & _T_1898; // @[Cache.scala 295:85]
  wire  _T_1900 = _T_1899 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_254 = _T_1900 | vArrayWire_28_0; // @[Reg.scala 28:19]
  wire  _T_1910 = selArrayWire_28 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1911 = _T_1894 & _T_1910; // @[Cache.scala 295:85]
  wire  _T_1912 = _T_1911 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_256 = _T_1912 | vArrayWire_28_1; // @[Reg.scala 28:19]
  wire  _T_1922 = selArrayWire_28 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1923 = _T_1894 & _T_1922; // @[Cache.scala 295:85]
  wire  _T_1924 = _T_1923 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_258 = _T_1924 | vArrayWire_28_2; // @[Reg.scala 28:19]
  wire  _T_1934 = selArrayWire_28 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1935 = _T_1894 & _T_1934; // @[Cache.scala 295:85]
  wire  _T_1936 = _T_1935 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_260 = _T_1936 | vArrayWire_28_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1945 = selArrayWire_29 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_1947 = io_cacheOut_r_last_i & _T_192; // @[Cache.scala 292:28]
  wire  _T_1951 = selArrayWire_29 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_1952 = _T_1947 & _T_1951; // @[Cache.scala 295:85]
  wire  _T_1953 = _T_1952 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_263 = _T_1953 | vArrayWire_29_0; // @[Reg.scala 28:19]
  wire  _T_1963 = selArrayWire_29 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_1964 = _T_1947 & _T_1963; // @[Cache.scala 295:85]
  wire  _T_1965 = _T_1964 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_265 = _T_1965 | vArrayWire_29_1; // @[Reg.scala 28:19]
  wire  _T_1975 = selArrayWire_29 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_1976 = _T_1947 & _T_1975; // @[Cache.scala 295:85]
  wire  _T_1977 = _T_1976 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_267 = _T_1977 | vArrayWire_29_2; // @[Reg.scala 28:19]
  wire  _T_1987 = selArrayWire_29 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_1988 = _T_1947 & _T_1987; // @[Cache.scala 295:85]
  wire  _T_1989 = _T_1988 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_269 = _T_1989 | vArrayWire_29_3; // @[Reg.scala 28:19]
  wire [1:0] _T_1998 = selArrayWire_30 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2000 = io_cacheOut_r_last_i & _T_194; // @[Cache.scala 292:28]
  wire  _T_2004 = selArrayWire_30 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2005 = _T_2000 & _T_2004; // @[Cache.scala 295:85]
  wire  _T_2006 = _T_2005 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_272 = _T_2006 | vArrayWire_30_0; // @[Reg.scala 28:19]
  wire  _T_2016 = selArrayWire_30 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2017 = _T_2000 & _T_2016; // @[Cache.scala 295:85]
  wire  _T_2018 = _T_2017 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_274 = _T_2018 | vArrayWire_30_1; // @[Reg.scala 28:19]
  wire  _T_2028 = selArrayWire_30 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2029 = _T_2000 & _T_2028; // @[Cache.scala 295:85]
  wire  _T_2030 = _T_2029 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_276 = _T_2030 | vArrayWire_30_2; // @[Reg.scala 28:19]
  wire  _T_2040 = selArrayWire_30 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2041 = _T_2000 & _T_2040; // @[Cache.scala 295:85]
  wire  _T_2042 = _T_2041 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_278 = _T_2042 | vArrayWire_30_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2051 = selArrayWire_31 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2053 = io_cacheOut_r_last_i & _T_196; // @[Cache.scala 292:28]
  wire  _T_2057 = selArrayWire_31 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2058 = _T_2053 & _T_2057; // @[Cache.scala 295:85]
  wire  _T_2059 = _T_2058 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_281 = _T_2059 | vArrayWire_31_0; // @[Reg.scala 28:19]
  wire  _T_2069 = selArrayWire_31 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2070 = _T_2053 & _T_2069; // @[Cache.scala 295:85]
  wire  _T_2071 = _T_2070 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_283 = _T_2071 | vArrayWire_31_1; // @[Reg.scala 28:19]
  wire  _T_2081 = selArrayWire_31 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2082 = _T_2053 & _T_2081; // @[Cache.scala 295:85]
  wire  _T_2083 = _T_2082 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_285 = _T_2083 | vArrayWire_31_2; // @[Reg.scala 28:19]
  wire  _T_2093 = selArrayWire_31 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2094 = _T_2053 & _T_2093; // @[Cache.scala 295:85]
  wire  _T_2095 = _T_2094 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_287 = _T_2095 | vArrayWire_31_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2104 = selArrayWire_32 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2106 = io_cacheOut_r_last_i & _T_198; // @[Cache.scala 292:28]
  wire  _T_2110 = selArrayWire_32 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2111 = _T_2106 & _T_2110; // @[Cache.scala 295:85]
  wire  _T_2112 = _T_2111 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_290 = _T_2112 | vArrayWire_32_0; // @[Reg.scala 28:19]
  wire  _T_2122 = selArrayWire_32 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2123 = _T_2106 & _T_2122; // @[Cache.scala 295:85]
  wire  _T_2124 = _T_2123 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_292 = _T_2124 | vArrayWire_32_1; // @[Reg.scala 28:19]
  wire  _T_2134 = selArrayWire_32 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2135 = _T_2106 & _T_2134; // @[Cache.scala 295:85]
  wire  _T_2136 = _T_2135 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_294 = _T_2136 | vArrayWire_32_2; // @[Reg.scala 28:19]
  wire  _T_2146 = selArrayWire_32 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2147 = _T_2106 & _T_2146; // @[Cache.scala 295:85]
  wire  _T_2148 = _T_2147 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_296 = _T_2148 | vArrayWire_32_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2157 = selArrayWire_33 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2159 = io_cacheOut_r_last_i & _T_200; // @[Cache.scala 292:28]
  wire  _T_2163 = selArrayWire_33 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2164 = _T_2159 & _T_2163; // @[Cache.scala 295:85]
  wire  _T_2165 = _T_2164 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_299 = _T_2165 | vArrayWire_33_0; // @[Reg.scala 28:19]
  wire  _T_2175 = selArrayWire_33 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2176 = _T_2159 & _T_2175; // @[Cache.scala 295:85]
  wire  _T_2177 = _T_2176 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_301 = _T_2177 | vArrayWire_33_1; // @[Reg.scala 28:19]
  wire  _T_2187 = selArrayWire_33 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2188 = _T_2159 & _T_2187; // @[Cache.scala 295:85]
  wire  _T_2189 = _T_2188 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_303 = _T_2189 | vArrayWire_33_2; // @[Reg.scala 28:19]
  wire  _T_2199 = selArrayWire_33 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2200 = _T_2159 & _T_2199; // @[Cache.scala 295:85]
  wire  _T_2201 = _T_2200 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_305 = _T_2201 | vArrayWire_33_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2210 = selArrayWire_34 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2212 = io_cacheOut_r_last_i & _T_202; // @[Cache.scala 292:28]
  wire  _T_2216 = selArrayWire_34 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2217 = _T_2212 & _T_2216; // @[Cache.scala 295:85]
  wire  _T_2218 = _T_2217 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_308 = _T_2218 | vArrayWire_34_0; // @[Reg.scala 28:19]
  wire  _T_2228 = selArrayWire_34 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2229 = _T_2212 & _T_2228; // @[Cache.scala 295:85]
  wire  _T_2230 = _T_2229 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_310 = _T_2230 | vArrayWire_34_1; // @[Reg.scala 28:19]
  wire  _T_2240 = selArrayWire_34 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2241 = _T_2212 & _T_2240; // @[Cache.scala 295:85]
  wire  _T_2242 = _T_2241 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_312 = _T_2242 | vArrayWire_34_2; // @[Reg.scala 28:19]
  wire  _T_2252 = selArrayWire_34 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2253 = _T_2212 & _T_2252; // @[Cache.scala 295:85]
  wire  _T_2254 = _T_2253 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_314 = _T_2254 | vArrayWire_34_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2263 = selArrayWire_35 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2265 = io_cacheOut_r_last_i & _T_204; // @[Cache.scala 292:28]
  wire  _T_2269 = selArrayWire_35 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2270 = _T_2265 & _T_2269; // @[Cache.scala 295:85]
  wire  _T_2271 = _T_2270 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_317 = _T_2271 | vArrayWire_35_0; // @[Reg.scala 28:19]
  wire  _T_2281 = selArrayWire_35 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2282 = _T_2265 & _T_2281; // @[Cache.scala 295:85]
  wire  _T_2283 = _T_2282 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_319 = _T_2283 | vArrayWire_35_1; // @[Reg.scala 28:19]
  wire  _T_2293 = selArrayWire_35 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2294 = _T_2265 & _T_2293; // @[Cache.scala 295:85]
  wire  _T_2295 = _T_2294 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_321 = _T_2295 | vArrayWire_35_2; // @[Reg.scala 28:19]
  wire  _T_2305 = selArrayWire_35 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2306 = _T_2265 & _T_2305; // @[Cache.scala 295:85]
  wire  _T_2307 = _T_2306 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_323 = _T_2307 | vArrayWire_35_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2316 = selArrayWire_36 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2318 = io_cacheOut_r_last_i & _T_206; // @[Cache.scala 292:28]
  wire  _T_2322 = selArrayWire_36 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2323 = _T_2318 & _T_2322; // @[Cache.scala 295:85]
  wire  _T_2324 = _T_2323 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_326 = _T_2324 | vArrayWire_36_0; // @[Reg.scala 28:19]
  wire  _T_2334 = selArrayWire_36 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2335 = _T_2318 & _T_2334; // @[Cache.scala 295:85]
  wire  _T_2336 = _T_2335 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_328 = _T_2336 | vArrayWire_36_1; // @[Reg.scala 28:19]
  wire  _T_2346 = selArrayWire_36 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2347 = _T_2318 & _T_2346; // @[Cache.scala 295:85]
  wire  _T_2348 = _T_2347 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_330 = _T_2348 | vArrayWire_36_2; // @[Reg.scala 28:19]
  wire  _T_2358 = selArrayWire_36 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2359 = _T_2318 & _T_2358; // @[Cache.scala 295:85]
  wire  _T_2360 = _T_2359 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_332 = _T_2360 | vArrayWire_36_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2369 = selArrayWire_37 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2371 = io_cacheOut_r_last_i & _T_208; // @[Cache.scala 292:28]
  wire  _T_2375 = selArrayWire_37 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2376 = _T_2371 & _T_2375; // @[Cache.scala 295:85]
  wire  _T_2377 = _T_2376 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_335 = _T_2377 | vArrayWire_37_0; // @[Reg.scala 28:19]
  wire  _T_2387 = selArrayWire_37 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2388 = _T_2371 & _T_2387; // @[Cache.scala 295:85]
  wire  _T_2389 = _T_2388 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_337 = _T_2389 | vArrayWire_37_1; // @[Reg.scala 28:19]
  wire  _T_2399 = selArrayWire_37 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2400 = _T_2371 & _T_2399; // @[Cache.scala 295:85]
  wire  _T_2401 = _T_2400 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_339 = _T_2401 | vArrayWire_37_2; // @[Reg.scala 28:19]
  wire  _T_2411 = selArrayWire_37 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2412 = _T_2371 & _T_2411; // @[Cache.scala 295:85]
  wire  _T_2413 = _T_2412 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_341 = _T_2413 | vArrayWire_37_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2422 = selArrayWire_38 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2424 = io_cacheOut_r_last_i & _T_210; // @[Cache.scala 292:28]
  wire  _T_2428 = selArrayWire_38 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2429 = _T_2424 & _T_2428; // @[Cache.scala 295:85]
  wire  _T_2430 = _T_2429 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_344 = _T_2430 | vArrayWire_38_0; // @[Reg.scala 28:19]
  wire  _T_2440 = selArrayWire_38 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2441 = _T_2424 & _T_2440; // @[Cache.scala 295:85]
  wire  _T_2442 = _T_2441 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_346 = _T_2442 | vArrayWire_38_1; // @[Reg.scala 28:19]
  wire  _T_2452 = selArrayWire_38 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2453 = _T_2424 & _T_2452; // @[Cache.scala 295:85]
  wire  _T_2454 = _T_2453 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_348 = _T_2454 | vArrayWire_38_2; // @[Reg.scala 28:19]
  wire  _T_2464 = selArrayWire_38 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2465 = _T_2424 & _T_2464; // @[Cache.scala 295:85]
  wire  _T_2466 = _T_2465 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_350 = _T_2466 | vArrayWire_38_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2475 = selArrayWire_39 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2477 = io_cacheOut_r_last_i & _T_212; // @[Cache.scala 292:28]
  wire  _T_2481 = selArrayWire_39 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2482 = _T_2477 & _T_2481; // @[Cache.scala 295:85]
  wire  _T_2483 = _T_2482 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_353 = _T_2483 | vArrayWire_39_0; // @[Reg.scala 28:19]
  wire  _T_2493 = selArrayWire_39 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2494 = _T_2477 & _T_2493; // @[Cache.scala 295:85]
  wire  _T_2495 = _T_2494 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_355 = _T_2495 | vArrayWire_39_1; // @[Reg.scala 28:19]
  wire  _T_2505 = selArrayWire_39 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2506 = _T_2477 & _T_2505; // @[Cache.scala 295:85]
  wire  _T_2507 = _T_2506 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_357 = _T_2507 | vArrayWire_39_2; // @[Reg.scala 28:19]
  wire  _T_2517 = selArrayWire_39 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2518 = _T_2477 & _T_2517; // @[Cache.scala 295:85]
  wire  _T_2519 = _T_2518 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_359 = _T_2519 | vArrayWire_39_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2528 = selArrayWire_40 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2530 = io_cacheOut_r_last_i & _T_214; // @[Cache.scala 292:28]
  wire  _T_2534 = selArrayWire_40 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2535 = _T_2530 & _T_2534; // @[Cache.scala 295:85]
  wire  _T_2536 = _T_2535 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_362 = _T_2536 | vArrayWire_40_0; // @[Reg.scala 28:19]
  wire  _T_2546 = selArrayWire_40 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2547 = _T_2530 & _T_2546; // @[Cache.scala 295:85]
  wire  _T_2548 = _T_2547 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_364 = _T_2548 | vArrayWire_40_1; // @[Reg.scala 28:19]
  wire  _T_2558 = selArrayWire_40 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2559 = _T_2530 & _T_2558; // @[Cache.scala 295:85]
  wire  _T_2560 = _T_2559 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_366 = _T_2560 | vArrayWire_40_2; // @[Reg.scala 28:19]
  wire  _T_2570 = selArrayWire_40 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2571 = _T_2530 & _T_2570; // @[Cache.scala 295:85]
  wire  _T_2572 = _T_2571 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_368 = _T_2572 | vArrayWire_40_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2581 = selArrayWire_41 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2583 = io_cacheOut_r_last_i & _T_216; // @[Cache.scala 292:28]
  wire  _T_2587 = selArrayWire_41 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2588 = _T_2583 & _T_2587; // @[Cache.scala 295:85]
  wire  _T_2589 = _T_2588 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_371 = _T_2589 | vArrayWire_41_0; // @[Reg.scala 28:19]
  wire  _T_2599 = selArrayWire_41 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2600 = _T_2583 & _T_2599; // @[Cache.scala 295:85]
  wire  _T_2601 = _T_2600 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_373 = _T_2601 | vArrayWire_41_1; // @[Reg.scala 28:19]
  wire  _T_2611 = selArrayWire_41 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2612 = _T_2583 & _T_2611; // @[Cache.scala 295:85]
  wire  _T_2613 = _T_2612 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_375 = _T_2613 | vArrayWire_41_2; // @[Reg.scala 28:19]
  wire  _T_2623 = selArrayWire_41 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2624 = _T_2583 & _T_2623; // @[Cache.scala 295:85]
  wire  _T_2625 = _T_2624 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_377 = _T_2625 | vArrayWire_41_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2634 = selArrayWire_42 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2636 = io_cacheOut_r_last_i & _T_218; // @[Cache.scala 292:28]
  wire  _T_2640 = selArrayWire_42 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2641 = _T_2636 & _T_2640; // @[Cache.scala 295:85]
  wire  _T_2642 = _T_2641 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_380 = _T_2642 | vArrayWire_42_0; // @[Reg.scala 28:19]
  wire  _T_2652 = selArrayWire_42 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2653 = _T_2636 & _T_2652; // @[Cache.scala 295:85]
  wire  _T_2654 = _T_2653 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_382 = _T_2654 | vArrayWire_42_1; // @[Reg.scala 28:19]
  wire  _T_2664 = selArrayWire_42 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2665 = _T_2636 & _T_2664; // @[Cache.scala 295:85]
  wire  _T_2666 = _T_2665 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_384 = _T_2666 | vArrayWire_42_2; // @[Reg.scala 28:19]
  wire  _T_2676 = selArrayWire_42 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2677 = _T_2636 & _T_2676; // @[Cache.scala 295:85]
  wire  _T_2678 = _T_2677 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_386 = _T_2678 | vArrayWire_42_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2687 = selArrayWire_43 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2689 = io_cacheOut_r_last_i & _T_220; // @[Cache.scala 292:28]
  wire  _T_2693 = selArrayWire_43 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2694 = _T_2689 & _T_2693; // @[Cache.scala 295:85]
  wire  _T_2695 = _T_2694 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_389 = _T_2695 | vArrayWire_43_0; // @[Reg.scala 28:19]
  wire  _T_2705 = selArrayWire_43 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2706 = _T_2689 & _T_2705; // @[Cache.scala 295:85]
  wire  _T_2707 = _T_2706 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_391 = _T_2707 | vArrayWire_43_1; // @[Reg.scala 28:19]
  wire  _T_2717 = selArrayWire_43 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2718 = _T_2689 & _T_2717; // @[Cache.scala 295:85]
  wire  _T_2719 = _T_2718 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_393 = _T_2719 | vArrayWire_43_2; // @[Reg.scala 28:19]
  wire  _T_2729 = selArrayWire_43 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2730 = _T_2689 & _T_2729; // @[Cache.scala 295:85]
  wire  _T_2731 = _T_2730 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_395 = _T_2731 | vArrayWire_43_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2740 = selArrayWire_44 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2742 = io_cacheOut_r_last_i & _T_222; // @[Cache.scala 292:28]
  wire  _T_2746 = selArrayWire_44 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2747 = _T_2742 & _T_2746; // @[Cache.scala 295:85]
  wire  _T_2748 = _T_2747 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_398 = _T_2748 | vArrayWire_44_0; // @[Reg.scala 28:19]
  wire  _T_2758 = selArrayWire_44 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2759 = _T_2742 & _T_2758; // @[Cache.scala 295:85]
  wire  _T_2760 = _T_2759 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_400 = _T_2760 | vArrayWire_44_1; // @[Reg.scala 28:19]
  wire  _T_2770 = selArrayWire_44 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2771 = _T_2742 & _T_2770; // @[Cache.scala 295:85]
  wire  _T_2772 = _T_2771 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_402 = _T_2772 | vArrayWire_44_2; // @[Reg.scala 28:19]
  wire  _T_2782 = selArrayWire_44 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2783 = _T_2742 & _T_2782; // @[Cache.scala 295:85]
  wire  _T_2784 = _T_2783 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_404 = _T_2784 | vArrayWire_44_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2793 = selArrayWire_45 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2795 = io_cacheOut_r_last_i & _T_224; // @[Cache.scala 292:28]
  wire  _T_2799 = selArrayWire_45 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2800 = _T_2795 & _T_2799; // @[Cache.scala 295:85]
  wire  _T_2801 = _T_2800 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_407 = _T_2801 | vArrayWire_45_0; // @[Reg.scala 28:19]
  wire  _T_2811 = selArrayWire_45 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2812 = _T_2795 & _T_2811; // @[Cache.scala 295:85]
  wire  _T_2813 = _T_2812 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_409 = _T_2813 | vArrayWire_45_1; // @[Reg.scala 28:19]
  wire  _T_2823 = selArrayWire_45 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2824 = _T_2795 & _T_2823; // @[Cache.scala 295:85]
  wire  _T_2825 = _T_2824 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_411 = _T_2825 | vArrayWire_45_2; // @[Reg.scala 28:19]
  wire  _T_2835 = selArrayWire_45 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2836 = _T_2795 & _T_2835; // @[Cache.scala 295:85]
  wire  _T_2837 = _T_2836 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_413 = _T_2837 | vArrayWire_45_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2846 = selArrayWire_46 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2848 = io_cacheOut_r_last_i & _T_226; // @[Cache.scala 292:28]
  wire  _T_2852 = selArrayWire_46 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2853 = _T_2848 & _T_2852; // @[Cache.scala 295:85]
  wire  _T_2854 = _T_2853 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_416 = _T_2854 | vArrayWire_46_0; // @[Reg.scala 28:19]
  wire  _T_2864 = selArrayWire_46 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2865 = _T_2848 & _T_2864; // @[Cache.scala 295:85]
  wire  _T_2866 = _T_2865 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_418 = _T_2866 | vArrayWire_46_1; // @[Reg.scala 28:19]
  wire  _T_2876 = selArrayWire_46 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2877 = _T_2848 & _T_2876; // @[Cache.scala 295:85]
  wire  _T_2878 = _T_2877 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_420 = _T_2878 | vArrayWire_46_2; // @[Reg.scala 28:19]
  wire  _T_2888 = selArrayWire_46 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2889 = _T_2848 & _T_2888; // @[Cache.scala 295:85]
  wire  _T_2890 = _T_2889 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_422 = _T_2890 | vArrayWire_46_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2899 = selArrayWire_47 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2901 = io_cacheOut_r_last_i & _T_228; // @[Cache.scala 292:28]
  wire  _T_2905 = selArrayWire_47 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2906 = _T_2901 & _T_2905; // @[Cache.scala 295:85]
  wire  _T_2907 = _T_2906 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_425 = _T_2907 | vArrayWire_47_0; // @[Reg.scala 28:19]
  wire  _T_2917 = selArrayWire_47 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2918 = _T_2901 & _T_2917; // @[Cache.scala 295:85]
  wire  _T_2919 = _T_2918 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_427 = _T_2919 | vArrayWire_47_1; // @[Reg.scala 28:19]
  wire  _T_2929 = selArrayWire_47 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2930 = _T_2901 & _T_2929; // @[Cache.scala 295:85]
  wire  _T_2931 = _T_2930 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_429 = _T_2931 | vArrayWire_47_2; // @[Reg.scala 28:19]
  wire  _T_2941 = selArrayWire_47 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2942 = _T_2901 & _T_2941; // @[Cache.scala 295:85]
  wire  _T_2943 = _T_2942 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_431 = _T_2943 | vArrayWire_47_3; // @[Reg.scala 28:19]
  wire [1:0] _T_2952 = selArrayWire_48 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_2954 = io_cacheOut_r_last_i & _T_230; // @[Cache.scala 292:28]
  wire  _T_2958 = selArrayWire_48 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_2959 = _T_2954 & _T_2958; // @[Cache.scala 295:85]
  wire  _T_2960 = _T_2959 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_434 = _T_2960 | vArrayWire_48_0; // @[Reg.scala 28:19]
  wire  _T_2970 = selArrayWire_48 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_2971 = _T_2954 & _T_2970; // @[Cache.scala 295:85]
  wire  _T_2972 = _T_2971 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_436 = _T_2972 | vArrayWire_48_1; // @[Reg.scala 28:19]
  wire  _T_2982 = selArrayWire_48 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_2983 = _T_2954 & _T_2982; // @[Cache.scala 295:85]
  wire  _T_2984 = _T_2983 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_438 = _T_2984 | vArrayWire_48_2; // @[Reg.scala 28:19]
  wire  _T_2994 = selArrayWire_48 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_2995 = _T_2954 & _T_2994; // @[Cache.scala 295:85]
  wire  _T_2996 = _T_2995 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_440 = _T_2996 | vArrayWire_48_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3005 = selArrayWire_49 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3007 = io_cacheOut_r_last_i & _T_232; // @[Cache.scala 292:28]
  wire  _T_3011 = selArrayWire_49 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3012 = _T_3007 & _T_3011; // @[Cache.scala 295:85]
  wire  _T_3013 = _T_3012 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_443 = _T_3013 | vArrayWire_49_0; // @[Reg.scala 28:19]
  wire  _T_3023 = selArrayWire_49 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3024 = _T_3007 & _T_3023; // @[Cache.scala 295:85]
  wire  _T_3025 = _T_3024 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_445 = _T_3025 | vArrayWire_49_1; // @[Reg.scala 28:19]
  wire  _T_3035 = selArrayWire_49 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3036 = _T_3007 & _T_3035; // @[Cache.scala 295:85]
  wire  _T_3037 = _T_3036 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_447 = _T_3037 | vArrayWire_49_2; // @[Reg.scala 28:19]
  wire  _T_3047 = selArrayWire_49 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3048 = _T_3007 & _T_3047; // @[Cache.scala 295:85]
  wire  _T_3049 = _T_3048 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_449 = _T_3049 | vArrayWire_49_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3058 = selArrayWire_50 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3060 = io_cacheOut_r_last_i & _T_234; // @[Cache.scala 292:28]
  wire  _T_3064 = selArrayWire_50 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3065 = _T_3060 & _T_3064; // @[Cache.scala 295:85]
  wire  _T_3066 = _T_3065 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_452 = _T_3066 | vArrayWire_50_0; // @[Reg.scala 28:19]
  wire  _T_3076 = selArrayWire_50 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3077 = _T_3060 & _T_3076; // @[Cache.scala 295:85]
  wire  _T_3078 = _T_3077 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_454 = _T_3078 | vArrayWire_50_1; // @[Reg.scala 28:19]
  wire  _T_3088 = selArrayWire_50 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3089 = _T_3060 & _T_3088; // @[Cache.scala 295:85]
  wire  _T_3090 = _T_3089 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_456 = _T_3090 | vArrayWire_50_2; // @[Reg.scala 28:19]
  wire  _T_3100 = selArrayWire_50 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3101 = _T_3060 & _T_3100; // @[Cache.scala 295:85]
  wire  _T_3102 = _T_3101 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_458 = _T_3102 | vArrayWire_50_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3111 = selArrayWire_51 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3113 = io_cacheOut_r_last_i & _T_236; // @[Cache.scala 292:28]
  wire  _T_3117 = selArrayWire_51 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3118 = _T_3113 & _T_3117; // @[Cache.scala 295:85]
  wire  _T_3119 = _T_3118 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_461 = _T_3119 | vArrayWire_51_0; // @[Reg.scala 28:19]
  wire  _T_3129 = selArrayWire_51 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3130 = _T_3113 & _T_3129; // @[Cache.scala 295:85]
  wire  _T_3131 = _T_3130 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_463 = _T_3131 | vArrayWire_51_1; // @[Reg.scala 28:19]
  wire  _T_3141 = selArrayWire_51 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3142 = _T_3113 & _T_3141; // @[Cache.scala 295:85]
  wire  _T_3143 = _T_3142 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_465 = _T_3143 | vArrayWire_51_2; // @[Reg.scala 28:19]
  wire  _T_3153 = selArrayWire_51 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3154 = _T_3113 & _T_3153; // @[Cache.scala 295:85]
  wire  _T_3155 = _T_3154 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_467 = _T_3155 | vArrayWire_51_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3164 = selArrayWire_52 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3166 = io_cacheOut_r_last_i & _T_238; // @[Cache.scala 292:28]
  wire  _T_3170 = selArrayWire_52 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3171 = _T_3166 & _T_3170; // @[Cache.scala 295:85]
  wire  _T_3172 = _T_3171 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_470 = _T_3172 | vArrayWire_52_0; // @[Reg.scala 28:19]
  wire  _T_3182 = selArrayWire_52 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3183 = _T_3166 & _T_3182; // @[Cache.scala 295:85]
  wire  _T_3184 = _T_3183 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_472 = _T_3184 | vArrayWire_52_1; // @[Reg.scala 28:19]
  wire  _T_3194 = selArrayWire_52 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3195 = _T_3166 & _T_3194; // @[Cache.scala 295:85]
  wire  _T_3196 = _T_3195 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_474 = _T_3196 | vArrayWire_52_2; // @[Reg.scala 28:19]
  wire  _T_3206 = selArrayWire_52 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3207 = _T_3166 & _T_3206; // @[Cache.scala 295:85]
  wire  _T_3208 = _T_3207 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_476 = _T_3208 | vArrayWire_52_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3217 = selArrayWire_53 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3219 = io_cacheOut_r_last_i & _T_240; // @[Cache.scala 292:28]
  wire  _T_3223 = selArrayWire_53 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3224 = _T_3219 & _T_3223; // @[Cache.scala 295:85]
  wire  _T_3225 = _T_3224 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_479 = _T_3225 | vArrayWire_53_0; // @[Reg.scala 28:19]
  wire  _T_3235 = selArrayWire_53 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3236 = _T_3219 & _T_3235; // @[Cache.scala 295:85]
  wire  _T_3237 = _T_3236 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_481 = _T_3237 | vArrayWire_53_1; // @[Reg.scala 28:19]
  wire  _T_3247 = selArrayWire_53 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3248 = _T_3219 & _T_3247; // @[Cache.scala 295:85]
  wire  _T_3249 = _T_3248 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_483 = _T_3249 | vArrayWire_53_2; // @[Reg.scala 28:19]
  wire  _T_3259 = selArrayWire_53 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3260 = _T_3219 & _T_3259; // @[Cache.scala 295:85]
  wire  _T_3261 = _T_3260 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_485 = _T_3261 | vArrayWire_53_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3270 = selArrayWire_54 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3272 = io_cacheOut_r_last_i & _T_242; // @[Cache.scala 292:28]
  wire  _T_3276 = selArrayWire_54 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3277 = _T_3272 & _T_3276; // @[Cache.scala 295:85]
  wire  _T_3278 = _T_3277 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_488 = _T_3278 | vArrayWire_54_0; // @[Reg.scala 28:19]
  wire  _T_3288 = selArrayWire_54 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3289 = _T_3272 & _T_3288; // @[Cache.scala 295:85]
  wire  _T_3290 = _T_3289 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_490 = _T_3290 | vArrayWire_54_1; // @[Reg.scala 28:19]
  wire  _T_3300 = selArrayWire_54 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3301 = _T_3272 & _T_3300; // @[Cache.scala 295:85]
  wire  _T_3302 = _T_3301 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_492 = _T_3302 | vArrayWire_54_2; // @[Reg.scala 28:19]
  wire  _T_3312 = selArrayWire_54 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3313 = _T_3272 & _T_3312; // @[Cache.scala 295:85]
  wire  _T_3314 = _T_3313 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_494 = _T_3314 | vArrayWire_54_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3323 = selArrayWire_55 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3325 = io_cacheOut_r_last_i & _T_244; // @[Cache.scala 292:28]
  wire  _T_3329 = selArrayWire_55 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3330 = _T_3325 & _T_3329; // @[Cache.scala 295:85]
  wire  _T_3331 = _T_3330 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_497 = _T_3331 | vArrayWire_55_0; // @[Reg.scala 28:19]
  wire  _T_3341 = selArrayWire_55 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3342 = _T_3325 & _T_3341; // @[Cache.scala 295:85]
  wire  _T_3343 = _T_3342 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_499 = _T_3343 | vArrayWire_55_1; // @[Reg.scala 28:19]
  wire  _T_3353 = selArrayWire_55 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3354 = _T_3325 & _T_3353; // @[Cache.scala 295:85]
  wire  _T_3355 = _T_3354 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_501 = _T_3355 | vArrayWire_55_2; // @[Reg.scala 28:19]
  wire  _T_3365 = selArrayWire_55 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3366 = _T_3325 & _T_3365; // @[Cache.scala 295:85]
  wire  _T_3367 = _T_3366 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_503 = _T_3367 | vArrayWire_55_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3376 = selArrayWire_56 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3378 = io_cacheOut_r_last_i & _T_246; // @[Cache.scala 292:28]
  wire  _T_3382 = selArrayWire_56 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3383 = _T_3378 & _T_3382; // @[Cache.scala 295:85]
  wire  _T_3384 = _T_3383 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_506 = _T_3384 | vArrayWire_56_0; // @[Reg.scala 28:19]
  wire  _T_3394 = selArrayWire_56 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3395 = _T_3378 & _T_3394; // @[Cache.scala 295:85]
  wire  _T_3396 = _T_3395 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_508 = _T_3396 | vArrayWire_56_1; // @[Reg.scala 28:19]
  wire  _T_3406 = selArrayWire_56 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3407 = _T_3378 & _T_3406; // @[Cache.scala 295:85]
  wire  _T_3408 = _T_3407 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_510 = _T_3408 | vArrayWire_56_2; // @[Reg.scala 28:19]
  wire  _T_3418 = selArrayWire_56 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3419 = _T_3378 & _T_3418; // @[Cache.scala 295:85]
  wire  _T_3420 = _T_3419 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_512 = _T_3420 | vArrayWire_56_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3429 = selArrayWire_57 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3431 = io_cacheOut_r_last_i & _T_248; // @[Cache.scala 292:28]
  wire  _T_3435 = selArrayWire_57 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3436 = _T_3431 & _T_3435; // @[Cache.scala 295:85]
  wire  _T_3437 = _T_3436 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_515 = _T_3437 | vArrayWire_57_0; // @[Reg.scala 28:19]
  wire  _T_3447 = selArrayWire_57 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3448 = _T_3431 & _T_3447; // @[Cache.scala 295:85]
  wire  _T_3449 = _T_3448 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_517 = _T_3449 | vArrayWire_57_1; // @[Reg.scala 28:19]
  wire  _T_3459 = selArrayWire_57 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3460 = _T_3431 & _T_3459; // @[Cache.scala 295:85]
  wire  _T_3461 = _T_3460 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_519 = _T_3461 | vArrayWire_57_2; // @[Reg.scala 28:19]
  wire  _T_3471 = selArrayWire_57 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3472 = _T_3431 & _T_3471; // @[Cache.scala 295:85]
  wire  _T_3473 = _T_3472 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_521 = _T_3473 | vArrayWire_57_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3482 = selArrayWire_58 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3484 = io_cacheOut_r_last_i & _T_250; // @[Cache.scala 292:28]
  wire  _T_3488 = selArrayWire_58 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3489 = _T_3484 & _T_3488; // @[Cache.scala 295:85]
  wire  _T_3490 = _T_3489 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_524 = _T_3490 | vArrayWire_58_0; // @[Reg.scala 28:19]
  wire  _T_3500 = selArrayWire_58 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3501 = _T_3484 & _T_3500; // @[Cache.scala 295:85]
  wire  _T_3502 = _T_3501 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_526 = _T_3502 | vArrayWire_58_1; // @[Reg.scala 28:19]
  wire  _T_3512 = selArrayWire_58 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3513 = _T_3484 & _T_3512; // @[Cache.scala 295:85]
  wire  _T_3514 = _T_3513 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_528 = _T_3514 | vArrayWire_58_2; // @[Reg.scala 28:19]
  wire  _T_3524 = selArrayWire_58 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3525 = _T_3484 & _T_3524; // @[Cache.scala 295:85]
  wire  _T_3526 = _T_3525 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_530 = _T_3526 | vArrayWire_58_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3535 = selArrayWire_59 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3537 = io_cacheOut_r_last_i & _T_252; // @[Cache.scala 292:28]
  wire  _T_3541 = selArrayWire_59 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3542 = _T_3537 & _T_3541; // @[Cache.scala 295:85]
  wire  _T_3543 = _T_3542 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_533 = _T_3543 | vArrayWire_59_0; // @[Reg.scala 28:19]
  wire  _T_3553 = selArrayWire_59 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3554 = _T_3537 & _T_3553; // @[Cache.scala 295:85]
  wire  _T_3555 = _T_3554 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_535 = _T_3555 | vArrayWire_59_1; // @[Reg.scala 28:19]
  wire  _T_3565 = selArrayWire_59 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3566 = _T_3537 & _T_3565; // @[Cache.scala 295:85]
  wire  _T_3567 = _T_3566 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_537 = _T_3567 | vArrayWire_59_2; // @[Reg.scala 28:19]
  wire  _T_3577 = selArrayWire_59 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3578 = _T_3537 & _T_3577; // @[Cache.scala 295:85]
  wire  _T_3579 = _T_3578 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_539 = _T_3579 | vArrayWire_59_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3588 = selArrayWire_60 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3590 = io_cacheOut_r_last_i & _T_254; // @[Cache.scala 292:28]
  wire  _T_3594 = selArrayWire_60 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3595 = _T_3590 & _T_3594; // @[Cache.scala 295:85]
  wire  _T_3596 = _T_3595 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_542 = _T_3596 | vArrayWire_60_0; // @[Reg.scala 28:19]
  wire  _T_3606 = selArrayWire_60 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3607 = _T_3590 & _T_3606; // @[Cache.scala 295:85]
  wire  _T_3608 = _T_3607 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_544 = _T_3608 | vArrayWire_60_1; // @[Reg.scala 28:19]
  wire  _T_3618 = selArrayWire_60 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3619 = _T_3590 & _T_3618; // @[Cache.scala 295:85]
  wire  _T_3620 = _T_3619 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_546 = _T_3620 | vArrayWire_60_2; // @[Reg.scala 28:19]
  wire  _T_3630 = selArrayWire_60 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3631 = _T_3590 & _T_3630; // @[Cache.scala 295:85]
  wire  _T_3632 = _T_3631 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_548 = _T_3632 | vArrayWire_60_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3641 = selArrayWire_61 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3643 = io_cacheOut_r_last_i & _T_256; // @[Cache.scala 292:28]
  wire  _T_3647 = selArrayWire_61 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3648 = _T_3643 & _T_3647; // @[Cache.scala 295:85]
  wire  _T_3649 = _T_3648 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_551 = _T_3649 | vArrayWire_61_0; // @[Reg.scala 28:19]
  wire  _T_3659 = selArrayWire_61 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3660 = _T_3643 & _T_3659; // @[Cache.scala 295:85]
  wire  _T_3661 = _T_3660 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_553 = _T_3661 | vArrayWire_61_1; // @[Reg.scala 28:19]
  wire  _T_3671 = selArrayWire_61 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3672 = _T_3643 & _T_3671; // @[Cache.scala 295:85]
  wire  _T_3673 = _T_3672 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_555 = _T_3673 | vArrayWire_61_2; // @[Reg.scala 28:19]
  wire  _T_3683 = selArrayWire_61 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3684 = _T_3643 & _T_3683; // @[Cache.scala 295:85]
  wire  _T_3685 = _T_3684 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_557 = _T_3685 | vArrayWire_61_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3694 = selArrayWire_62 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3696 = io_cacheOut_r_last_i & _T_258; // @[Cache.scala 292:28]
  wire  _T_3700 = selArrayWire_62 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3701 = _T_3696 & _T_3700; // @[Cache.scala 295:85]
  wire  _T_3702 = _T_3701 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_560 = _T_3702 | vArrayWire_62_0; // @[Reg.scala 28:19]
  wire  _T_3712 = selArrayWire_62 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3713 = _T_3696 & _T_3712; // @[Cache.scala 295:85]
  wire  _T_3714 = _T_3713 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_562 = _T_3714 | vArrayWire_62_1; // @[Reg.scala 28:19]
  wire  _T_3724 = selArrayWire_62 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3725 = _T_3696 & _T_3724; // @[Cache.scala 295:85]
  wire  _T_3726 = _T_3725 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_564 = _T_3726 | vArrayWire_62_2; // @[Reg.scala 28:19]
  wire  _T_3736 = selArrayWire_62 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3737 = _T_3696 & _T_3736; // @[Cache.scala 295:85]
  wire  _T_3738 = _T_3737 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_566 = _T_3738 | vArrayWire_62_3; // @[Reg.scala 28:19]
  wire [1:0] _T_3747 = selArrayWire_63 + 2'h1; // @[Cache.scala 290:23]
  wire  _T_3749 = io_cacheOut_r_last_i & _T_260; // @[Cache.scala 292:28]
  wire  _T_3753 = selArrayWire_63 == 2'h0; // @[Cache.scala 295:104]
  wire  _T_3754 = _T_3749 & _T_3753; // @[Cache.scala 295:85]
  wire  _T_3755 = _T_3754 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_569 = _T_3755 | vArrayWire_63_0; // @[Reg.scala 28:19]
  wire  _T_3765 = selArrayWire_63 == 2'h1; // @[Cache.scala 295:104]
  wire  _T_3766 = _T_3749 & _T_3765; // @[Cache.scala 295:85]
  wire  _T_3767 = _T_3766 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_571 = _T_3767 | vArrayWire_63_1; // @[Reg.scala 28:19]
  wire  _T_3777 = selArrayWire_63 == 2'h2; // @[Cache.scala 295:104]
  wire  _T_3778 = _T_3749 & _T_3777; // @[Cache.scala 295:85]
  wire  _T_3779 = _T_3778 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_573 = _T_3779 | vArrayWire_63_2; // @[Reg.scala 28:19]
  wire  _T_3789 = selArrayWire_63 == 2'h3; // @[Cache.scala 295:104]
  wire  _T_3790 = _T_3749 & _T_3789; // @[Cache.scala 295:85]
  wire  _T_3791 = _T_3790 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_575 = _T_3791 | vArrayWire_63_3; // @[Reg.scala 28:19]
  wire [7:0] maskWrite_0 = io_cacheIn_mask[0] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_1 = io_cacheIn_mask[1] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_2 = io_cacheIn_mask[2] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_3 = io_cacheIn_mask[3] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_4 = io_cacheIn_mask[4] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_5 = io_cacheIn_mask[5] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_6 = io_cacheIn_mask[6] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_7 = io_cacheIn_mask[7] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [127:0] _T_3841 = {maskWrite_7,maskWrite_6,maskWrite_5,maskWrite_4,maskWrite_3,maskWrite_2,maskWrite_1,maskWrite_0,64'hffffffffffffffff}; // @[Cat.scala 29:58]
  wire [127:0] _T_3851 = {64'hffffffffffffffff,maskWrite_7,maskWrite_6,maskWrite_5,maskWrite_4,maskWrite_3,maskWrite_2,maskWrite_1,maskWrite_0}; // @[Cat.scala 29:58]
  wire [127:0] ramMaskWrite = offset[3] ? _T_3841 : _T_3851; // @[Cache.scala 313:25]
  wire  _T_3854 = _T_1 & io_cacheIn_wen; // @[Cache.scala 331:59]
  wire  _T_3856 = io_cacheIn_valid & hitArray_0; // @[Cache.scala 341:36]
  wire  _T_3857 = _T_3856 & isIdle; // @[Cache.scala 341:53]
  wire  _T_3858 = isMiss & io_cacheOut_r_valid_i; // @[Cache.scala 341:76]
  wire  _T_3859 = 2'h0 == sramSel; // @[Cache.scala 341:111]
  wire  _T_3860 = _T_3858 & _T_3859; // @[Cache.scala 341:102]
  wire  _T_3861 = _T_3857 | _T_3860; // @[Cache.scala 341:64]
  wire  _T_3863 = io_cacheIn_wen & isIdle; // @[Cache.scala 343:34]
  wire  _T_3867 = _T_3863 | _T_3860; // @[Cache.scala 343:45]
  wire [127:0] _T_3869 = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_3870 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 29:58]
  wire [127:0] _T_3871 = io_cacheOut_r_last_i ? _T_3869 : _T_3870; // @[Cache.scala 346:10]
  wire [127:0] _T_3873 = {io_cacheIn_data_write,64'h0}; // @[Cat.scala 29:58]
  wire [127:0] _T_3874 = {64'h0,io_cacheIn_data_write}; // @[Cat.scala 29:58]
  wire [127:0] _T_3875 = offset[3] ? _T_3873 : _T_3874; // @[Cache.scala 347:10]
  wire [127:0] _T_3883 = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 351:10]
  wire  _T_3885 = io_cacheIn_valid & hitArray_1; // @[Cache.scala 341:36]
  wire  _T_3886 = _T_3885 & isIdle; // @[Cache.scala 341:53]
  wire  _T_3888 = 2'h1 == sramSel; // @[Cache.scala 341:111]
  wire  _T_3889 = _T_3858 & _T_3888; // @[Cache.scala 341:102]
  wire  _T_3890 = _T_3886 | _T_3889; // @[Cache.scala 341:64]
  wire  _T_3896 = _T_3863 | _T_3889; // @[Cache.scala 343:45]
  wire  _T_3914 = io_cacheIn_valid & hitArray_2; // @[Cache.scala 341:36]
  wire  _T_3915 = _T_3914 & isIdle; // @[Cache.scala 341:53]
  wire  _T_3917 = 2'h2 == sramSel; // @[Cache.scala 341:111]
  wire  _T_3918 = _T_3858 & _T_3917; // @[Cache.scala 341:102]
  wire  _T_3919 = _T_3915 | _T_3918; // @[Cache.scala 341:64]
  wire  _T_3925 = _T_3863 | _T_3918; // @[Cache.scala 343:45]
  wire  _T_3943 = io_cacheIn_valid & hitArray_3; // @[Cache.scala 341:36]
  wire  _T_3944 = _T_3943 & isIdle; // @[Cache.scala 341:53]
  wire  _T_3946 = 2'h3 == sramSel; // @[Cache.scala 341:111]
  wire  _T_3947 = _T_3858 & _T_3946; // @[Cache.scala 341:102]
  wire  _T_3948 = _T_3944 | _T_3947; // @[Cache.scala 341:64]
  wire  _T_3954 = _T_3863 | _T_3947; // @[Cache.scala 343:45]
  wire  _T_3972 = isWrite & io_cacheOut_w_ready_i; // @[Cache.scala 357:31]
  wire  _T_3973 = _T_3972 | isBlock; // @[Cache.scala 357:57]
  wire  _T_3974 = isIdle & hit; // @[Cache.scala 357:77]
  wire  _T_3975 = ~io_cacheIn_wen; // @[Cache.scala 357:86]
  wire  _T_3976 = _T_3974 & _T_3975; // @[Cache.scala 357:83]
  assign io_cacheOut_ar_valid_o = cacheState == 2'h1; // @[Cache.scala 276:26]
  assign io_cacheOut_ar_addr_o = {io_cacheIn_addr[31:4],4'h0}; // @[Cache.scala 275:25]
  assign io_cacheOut_ar_len_o = {{7'd0}, isMiss}; // @[Cache.scala 274:24]
  assign io_cacheOut_w_valid_o = _T_3854 & isIdle; // @[Cache.scala 331:25]
  assign io_cacheOut_w_data_o = io_cacheIn_data_write; // @[Cache.scala 332:24]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 333:24]
  assign io_cacheOut_w_mask_o = io_cacheIn_mask; // @[Cache.scala 334:24]
  assign io_cacheOut_wsize = io_cacheIn_rsize; // @[Cache.scala 359:21]
  assign io_cacheIn_ready = _T_3973 | _T_3976; // @[Cache.scala 357:20]
  assign io_cacheIn_data_read = offset[3] ? waysel[127:64] : waysel[63:0]; // @[Cache.scala 263:24]
  assign io_SRAMIO_0_cen = ~_T_3861; // @[Cache.scala 341:13]
  assign io_SRAMIO_0_wen = ~_T_3867; // @[Cache.scala 343:13]
  assign io_SRAMIO_0_wdata = isMiss ? _T_3871 : _T_3875; // @[Cache.scala 344:15]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 342:14]
  assign io_SRAMIO_0_wmask = isMiss ? _T_3883 : ramMaskWrite; // @[Cache.scala 349:15]
  assign io_SRAMIO_1_cen = ~_T_3890; // @[Cache.scala 341:13]
  assign io_SRAMIO_1_wen = ~_T_3896; // @[Cache.scala 343:13]
  assign io_SRAMIO_1_wdata = isMiss ? _T_3871 : _T_3875; // @[Cache.scala 344:15]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 342:14]
  assign io_SRAMIO_1_wmask = isMiss ? _T_3883 : ramMaskWrite; // @[Cache.scala 349:15]
  assign io_SRAMIO_2_cen = ~_T_3919; // @[Cache.scala 341:13]
  assign io_SRAMIO_2_wen = ~_T_3925; // @[Cache.scala 343:13]
  assign io_SRAMIO_2_wdata = isMiss ? _T_3871 : _T_3875; // @[Cache.scala 344:15]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 342:14]
  assign io_SRAMIO_2_wmask = isMiss ? _T_3883 : ramMaskWrite; // @[Cache.scala 349:15]
  assign io_SRAMIO_3_cen = ~_T_3948; // @[Cache.scala 341:13]
  assign io_SRAMIO_3_wen = ~_T_3954; // @[Cache.scala 343:13]
  assign io_SRAMIO_3_wdata = isMiss ? _T_3871 : _T_3875; // @[Cache.scala 344:15]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 342:14]
  assign io_SRAMIO_3_wmask = isMiss ? _T_3883 : ramMaskWrite; // @[Cache.scala 349:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cacheState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  vArrayWire_63_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vArrayWire_62_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  vArrayWire_61_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  vArrayWire_60_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vArrayWire_59_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  vArrayWire_58_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  vArrayWire_57_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  vArrayWire_56_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  vArrayWire_55_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  vArrayWire_54_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vArrayWire_53_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  vArrayWire_52_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  vArrayWire_51_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  vArrayWire_50_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  vArrayWire_49_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  vArrayWire_48_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  vArrayWire_47_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  vArrayWire_46_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  vArrayWire_45_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  vArrayWire_44_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  vArrayWire_43_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  vArrayWire_42_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  vArrayWire_41_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  vArrayWire_40_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  vArrayWire_39_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  vArrayWire_38_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vArrayWire_37_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  vArrayWire_36_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  vArrayWire_35_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  vArrayWire_34_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  vArrayWire_33_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  vArrayWire_32_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  vArrayWire_31_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  vArrayWire_30_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  vArrayWire_29_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  vArrayWire_28_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  vArrayWire_27_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  vArrayWire_26_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  vArrayWire_25_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  vArrayWire_24_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  vArrayWire_23_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  vArrayWire_22_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  vArrayWire_21_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  vArrayWire_20_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  vArrayWire_19_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  vArrayWire_18_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  vArrayWire_17_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  vArrayWire_16_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  vArrayWire_15_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  vArrayWire_14_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  vArrayWire_13_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  vArrayWire_12_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vArrayWire_11_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  vArrayWire_10_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  vArrayWire_9_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  vArrayWire_8_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  vArrayWire_7_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  vArrayWire_6_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  vArrayWire_5_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  vArrayWire_4_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  vArrayWire_3_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  vArrayWire_2_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  vArrayWire_1_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  vArrayWire_0_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tagArrayWire_63_0 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tagArrayWire_62_0 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tagArrayWire_61_0 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tagArrayWire_60_0 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tagArrayWire_59_0 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tagArrayWire_58_0 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tagArrayWire_57_0 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tagArrayWire_56_0 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tagArrayWire_55_0 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tagArrayWire_54_0 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tagArrayWire_53_0 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tagArrayWire_52_0 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tagArrayWire_51_0 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tagArrayWire_50_0 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tagArrayWire_49_0 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tagArrayWire_48_0 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tagArrayWire_47_0 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tagArrayWire_46_0 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tagArrayWire_45_0 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tagArrayWire_44_0 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tagArrayWire_43_0 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tagArrayWire_42_0 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tagArrayWire_41_0 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tagArrayWire_40_0 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tagArrayWire_39_0 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tagArrayWire_38_0 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tagArrayWire_37_0 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tagArrayWire_36_0 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tagArrayWire_35_0 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tagArrayWire_34_0 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tagArrayWire_33_0 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tagArrayWire_32_0 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tagArrayWire_31_0 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tagArrayWire_30_0 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tagArrayWire_29_0 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tagArrayWire_28_0 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tagArrayWire_27_0 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tagArrayWire_26_0 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tagArrayWire_25_0 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tagArrayWire_24_0 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tagArrayWire_23_0 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tagArrayWire_22_0 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tagArrayWire_21_0 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tagArrayWire_20_0 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tagArrayWire_19_0 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tagArrayWire_18_0 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tagArrayWire_17_0 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tagArrayWire_16_0 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tagArrayWire_15_0 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tagArrayWire_14_0 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tagArrayWire_13_0 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tagArrayWire_12_0 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tagArrayWire_11_0 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tagArrayWire_10_0 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tagArrayWire_9_0 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tagArrayWire_8_0 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tagArrayWire_7_0 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tagArrayWire_6_0 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tagArrayWire_5_0 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tagArrayWire_4_0 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tagArrayWire_3_0 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tagArrayWire_2_0 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tagArrayWire_1_0 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  tagArrayWire_0_0 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  vArrayWire_63_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  vArrayWire_62_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  vArrayWire_61_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  vArrayWire_60_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  vArrayWire_59_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  vArrayWire_58_1 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  vArrayWire_57_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  vArrayWire_56_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  vArrayWire_55_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  vArrayWire_54_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  vArrayWire_53_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  vArrayWire_52_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  vArrayWire_51_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  vArrayWire_50_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  vArrayWire_49_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  vArrayWire_48_1 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  vArrayWire_47_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  vArrayWire_46_1 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  vArrayWire_45_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  vArrayWire_44_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  vArrayWire_43_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  vArrayWire_42_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  vArrayWire_41_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  vArrayWire_40_1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  vArrayWire_39_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  vArrayWire_38_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  vArrayWire_37_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  vArrayWire_36_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  vArrayWire_35_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  vArrayWire_34_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  vArrayWire_33_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  vArrayWire_32_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  vArrayWire_31_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  vArrayWire_30_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  vArrayWire_29_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  vArrayWire_28_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  vArrayWire_27_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  vArrayWire_26_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  vArrayWire_25_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  vArrayWire_24_1 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  vArrayWire_23_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  vArrayWire_22_1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  vArrayWire_21_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  vArrayWire_20_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  vArrayWire_19_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  vArrayWire_18_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  vArrayWire_17_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  vArrayWire_16_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  vArrayWire_15_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  vArrayWire_14_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  vArrayWire_13_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  vArrayWire_12_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  vArrayWire_11_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  vArrayWire_10_1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vArrayWire_9_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  vArrayWire_8_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  vArrayWire_7_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  vArrayWire_6_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  vArrayWire_5_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  vArrayWire_4_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  vArrayWire_3_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  vArrayWire_2_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  vArrayWire_1_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  vArrayWire_0_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tagArrayWire_63_1 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  tagArrayWire_62_1 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  tagArrayWire_61_1 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  tagArrayWire_60_1 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  tagArrayWire_59_1 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  tagArrayWire_58_1 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  tagArrayWire_57_1 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  tagArrayWire_56_1 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  tagArrayWire_55_1 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  tagArrayWire_54_1 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  tagArrayWire_53_1 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  tagArrayWire_52_1 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  tagArrayWire_51_1 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  tagArrayWire_50_1 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  tagArrayWire_49_1 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  tagArrayWire_48_1 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  tagArrayWire_47_1 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  tagArrayWire_46_1 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  tagArrayWire_45_1 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  tagArrayWire_44_1 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  tagArrayWire_43_1 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  tagArrayWire_42_1 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  tagArrayWire_41_1 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  tagArrayWire_40_1 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  tagArrayWire_39_1 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  tagArrayWire_38_1 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  tagArrayWire_37_1 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  tagArrayWire_36_1 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  tagArrayWire_35_1 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  tagArrayWire_34_1 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  tagArrayWire_33_1 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  tagArrayWire_32_1 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  tagArrayWire_31_1 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  tagArrayWire_30_1 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  tagArrayWire_29_1 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  tagArrayWire_28_1 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  tagArrayWire_27_1 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  tagArrayWire_26_1 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  tagArrayWire_25_1 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  tagArrayWire_24_1 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  tagArrayWire_23_1 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  tagArrayWire_22_1 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  tagArrayWire_21_1 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  tagArrayWire_20_1 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  tagArrayWire_19_1 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  tagArrayWire_18_1 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  tagArrayWire_17_1 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  tagArrayWire_16_1 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  tagArrayWire_15_1 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  tagArrayWire_14_1 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  tagArrayWire_13_1 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  tagArrayWire_12_1 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  tagArrayWire_11_1 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  tagArrayWire_10_1 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  tagArrayWire_9_1 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  tagArrayWire_8_1 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  tagArrayWire_7_1 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  tagArrayWire_6_1 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  tagArrayWire_5_1 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  tagArrayWire_4_1 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  tagArrayWire_3_1 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  tagArrayWire_2_1 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  tagArrayWire_1_1 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  tagArrayWire_0_1 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  vArrayWire_63_2 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  vArrayWire_62_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  vArrayWire_61_2 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  vArrayWire_60_2 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  vArrayWire_59_2 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  vArrayWire_58_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  vArrayWire_57_2 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  vArrayWire_56_2 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  vArrayWire_55_2 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  vArrayWire_54_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  vArrayWire_53_2 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  vArrayWire_52_2 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  vArrayWire_51_2 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  vArrayWire_50_2 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  vArrayWire_49_2 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  vArrayWire_48_2 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  vArrayWire_47_2 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  vArrayWire_46_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  vArrayWire_45_2 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  vArrayWire_44_2 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  vArrayWire_43_2 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  vArrayWire_42_2 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  vArrayWire_41_2 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  vArrayWire_40_2 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  vArrayWire_39_2 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  vArrayWire_38_2 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  vArrayWire_37_2 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  vArrayWire_36_2 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  vArrayWire_35_2 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  vArrayWire_34_2 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  vArrayWire_33_2 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  vArrayWire_32_2 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  vArrayWire_31_2 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  vArrayWire_30_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  vArrayWire_29_2 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  vArrayWire_28_2 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  vArrayWire_27_2 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  vArrayWire_26_2 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  vArrayWire_25_2 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  vArrayWire_24_2 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  vArrayWire_23_2 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  vArrayWire_22_2 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  vArrayWire_21_2 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  vArrayWire_20_2 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  vArrayWire_19_2 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  vArrayWire_18_2 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  vArrayWire_17_2 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  vArrayWire_16_2 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  vArrayWire_15_2 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  vArrayWire_14_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  vArrayWire_13_2 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  vArrayWire_12_2 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  vArrayWire_11_2 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  vArrayWire_10_2 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  vArrayWire_9_2 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  vArrayWire_8_2 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  vArrayWire_7_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  vArrayWire_6_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  vArrayWire_5_2 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  vArrayWire_4_2 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  vArrayWire_3_2 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  vArrayWire_2_2 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  vArrayWire_1_2 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  vArrayWire_0_2 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  tagArrayWire_63_2 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  tagArrayWire_62_2 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  tagArrayWire_61_2 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  tagArrayWire_60_2 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  tagArrayWire_59_2 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  tagArrayWire_58_2 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  tagArrayWire_57_2 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  tagArrayWire_56_2 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  tagArrayWire_55_2 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  tagArrayWire_54_2 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  tagArrayWire_53_2 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  tagArrayWire_52_2 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  tagArrayWire_51_2 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  tagArrayWire_50_2 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  tagArrayWire_49_2 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  tagArrayWire_48_2 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  tagArrayWire_47_2 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  tagArrayWire_46_2 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  tagArrayWire_45_2 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  tagArrayWire_44_2 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  tagArrayWire_43_2 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  tagArrayWire_42_2 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  tagArrayWire_41_2 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  tagArrayWire_40_2 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  tagArrayWire_39_2 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  tagArrayWire_38_2 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  tagArrayWire_37_2 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  tagArrayWire_36_2 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  tagArrayWire_35_2 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  tagArrayWire_34_2 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  tagArrayWire_33_2 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  tagArrayWire_32_2 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  tagArrayWire_31_2 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  tagArrayWire_30_2 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  tagArrayWire_29_2 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  tagArrayWire_28_2 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  tagArrayWire_27_2 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  tagArrayWire_26_2 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  tagArrayWire_25_2 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  tagArrayWire_24_2 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  tagArrayWire_23_2 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  tagArrayWire_22_2 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  tagArrayWire_21_2 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  tagArrayWire_20_2 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  tagArrayWire_19_2 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  tagArrayWire_18_2 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  tagArrayWire_17_2 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  tagArrayWire_16_2 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  tagArrayWire_15_2 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  tagArrayWire_14_2 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  tagArrayWire_13_2 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  tagArrayWire_12_2 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  tagArrayWire_11_2 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  tagArrayWire_10_2 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  tagArrayWire_9_2 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  tagArrayWire_8_2 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  tagArrayWire_7_2 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  tagArrayWire_6_2 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  tagArrayWire_5_2 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  tagArrayWire_4_2 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  tagArrayWire_3_2 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  tagArrayWire_2_2 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  tagArrayWire_1_2 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  tagArrayWire_0_2 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  vArrayWire_63_3 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  vArrayWire_62_3 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  vArrayWire_61_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  vArrayWire_60_3 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  vArrayWire_59_3 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  vArrayWire_58_3 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  vArrayWire_57_3 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  vArrayWire_56_3 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  vArrayWire_55_3 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  vArrayWire_54_3 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  vArrayWire_53_3 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  vArrayWire_52_3 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  vArrayWire_51_3 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  vArrayWire_50_3 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  vArrayWire_49_3 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  vArrayWire_48_3 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  vArrayWire_47_3 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  vArrayWire_46_3 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  vArrayWire_45_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  vArrayWire_44_3 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  vArrayWire_43_3 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  vArrayWire_42_3 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  vArrayWire_41_3 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  vArrayWire_40_3 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  vArrayWire_39_3 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  vArrayWire_38_3 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  vArrayWire_37_3 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  vArrayWire_36_3 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  vArrayWire_35_3 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  vArrayWire_34_3 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  vArrayWire_33_3 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  vArrayWire_32_3 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  vArrayWire_31_3 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  vArrayWire_30_3 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  vArrayWire_29_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  vArrayWire_28_3 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  vArrayWire_27_3 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  vArrayWire_26_3 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  vArrayWire_25_3 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  vArrayWire_24_3 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  vArrayWire_23_3 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  vArrayWire_22_3 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  vArrayWire_21_3 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  vArrayWire_20_3 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  vArrayWire_19_3 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  vArrayWire_18_3 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  vArrayWire_17_3 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  vArrayWire_16_3 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  vArrayWire_15_3 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  vArrayWire_14_3 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  vArrayWire_13_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  vArrayWire_12_3 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  vArrayWire_11_3 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  vArrayWire_10_3 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  vArrayWire_9_3 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  vArrayWire_8_3 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  vArrayWire_7_3 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  vArrayWire_6_3 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  vArrayWire_5_3 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  vArrayWire_4_3 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  vArrayWire_3_3 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  vArrayWire_2_3 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  vArrayWire_1_3 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  vArrayWire_0_3 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  tagArrayWire_63_3 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  tagArrayWire_62_3 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  tagArrayWire_61_3 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  tagArrayWire_60_3 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  tagArrayWire_59_3 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  tagArrayWire_58_3 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  tagArrayWire_57_3 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  tagArrayWire_56_3 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  tagArrayWire_55_3 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  tagArrayWire_54_3 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  tagArrayWire_53_3 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  tagArrayWire_52_3 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  tagArrayWire_51_3 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  tagArrayWire_50_3 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  tagArrayWire_49_3 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  tagArrayWire_48_3 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  tagArrayWire_47_3 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  tagArrayWire_46_3 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  tagArrayWire_45_3 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  tagArrayWire_44_3 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  tagArrayWire_43_3 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  tagArrayWire_42_3 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  tagArrayWire_41_3 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  tagArrayWire_40_3 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  tagArrayWire_39_3 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  tagArrayWire_38_3 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  tagArrayWire_37_3 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  tagArrayWire_36_3 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  tagArrayWire_35_3 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  tagArrayWire_34_3 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  tagArrayWire_33_3 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  tagArrayWire_32_3 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  tagArrayWire_31_3 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  tagArrayWire_30_3 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  tagArrayWire_29_3 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  tagArrayWire_28_3 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  tagArrayWire_27_3 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  tagArrayWire_26_3 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  tagArrayWire_25_3 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  tagArrayWire_24_3 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  tagArrayWire_23_3 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  tagArrayWire_22_3 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  tagArrayWire_21_3 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  tagArrayWire_20_3 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  tagArrayWire_19_3 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  tagArrayWire_18_3 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  tagArrayWire_17_3 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  tagArrayWire_16_3 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  tagArrayWire_15_3 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  tagArrayWire_14_3 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  tagArrayWire_13_3 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  tagArrayWire_12_3 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  tagArrayWire_11_3 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  tagArrayWire_10_3 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  tagArrayWire_9_3 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  tagArrayWire_8_3 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  tagArrayWire_7_3 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  tagArrayWire_6_3 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  tagArrayWire_5_3 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  tagArrayWire_4_3 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  tagArrayWire_3_3 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  tagArrayWire_2_3 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  tagArrayWire_1_3 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  tagArrayWire_0_3 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  selArrayWire_1 = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  selArrayWire_0 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  selArrayWire_2 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  selArrayWire_3 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  selArrayWire_4 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  selArrayWire_5 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  selArrayWire_6 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  selArrayWire_7 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  selArrayWire_8 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  selArrayWire_9 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  selArrayWire_10 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  selArrayWire_11 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  selArrayWire_12 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  selArrayWire_13 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  selArrayWire_14 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  selArrayWire_15 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  selArrayWire_16 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  selArrayWire_17 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  selArrayWire_18 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  selArrayWire_19 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  selArrayWire_20 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  selArrayWire_21 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  selArrayWire_22 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  selArrayWire_23 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  selArrayWire_24 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  selArrayWire_25 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  selArrayWire_26 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  selArrayWire_27 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  selArrayWire_28 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  selArrayWire_29 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  selArrayWire_30 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  selArrayWire_31 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  selArrayWire_32 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  selArrayWire_33 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  selArrayWire_34 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  selArrayWire_35 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  selArrayWire_36 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  selArrayWire_37 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  selArrayWire_38 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  selArrayWire_39 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  selArrayWire_40 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  selArrayWire_41 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  selArrayWire_42 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  selArrayWire_43 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  selArrayWire_44 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  selArrayWire_45 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  selArrayWire_46 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  selArrayWire_47 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  selArrayWire_48 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  selArrayWire_49 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  selArrayWire_50 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  selArrayWire_51 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  selArrayWire_52 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  selArrayWire_53 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  selArrayWire_54 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  selArrayWire_55 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  selArrayWire_56 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  selArrayWire_57 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  selArrayWire_58 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  selArrayWire_59 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  selArrayWire_60 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  selArrayWire_61 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  selArrayWire_62 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  selArrayWire_63 = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cacheState <= 2'h0;
    end else if (_T_9) begin
      if (io_block) begin
        cacheState <= 2'h3;
      end else begin
        cacheState <= 2'h0;
      end
    end else if (_T_7) begin
      if (io_cacheOut_w_ready_i) begin
        if (io_block) begin
          cacheState <= 2'h3;
        end else begin
          cacheState <= 2'h0;
        end
      end else begin
        cacheState <= 2'h2;
      end
    end else if (_T_5) begin
      if (io_cacheOut_r_last_i) begin
        cacheState <= 2'h0;
      end else begin
        cacheState <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_cacheIn_wen) begin
        cacheState <= 2'h2;
      end else if (hit) begin
        cacheState <= 2'h0;
      end else begin
        cacheState <= 2'h1;
      end
    end else begin
      cacheState <= 2'h0;
    end
    if (reset) begin
      vArrayWire_63_0 <= 1'h0;
    end else begin
      vArrayWire_63_0 <= _GEN_569;
    end
    if (reset) begin
      vArrayWire_62_0 <= 1'h0;
    end else begin
      vArrayWire_62_0 <= _GEN_560;
    end
    if (reset) begin
      vArrayWire_61_0 <= 1'h0;
    end else begin
      vArrayWire_61_0 <= _GEN_551;
    end
    if (reset) begin
      vArrayWire_60_0 <= 1'h0;
    end else begin
      vArrayWire_60_0 <= _GEN_542;
    end
    if (reset) begin
      vArrayWire_59_0 <= 1'h0;
    end else begin
      vArrayWire_59_0 <= _GEN_533;
    end
    if (reset) begin
      vArrayWire_58_0 <= 1'h0;
    end else begin
      vArrayWire_58_0 <= _GEN_524;
    end
    if (reset) begin
      vArrayWire_57_0 <= 1'h0;
    end else begin
      vArrayWire_57_0 <= _GEN_515;
    end
    if (reset) begin
      vArrayWire_56_0 <= 1'h0;
    end else begin
      vArrayWire_56_0 <= _GEN_506;
    end
    if (reset) begin
      vArrayWire_55_0 <= 1'h0;
    end else begin
      vArrayWire_55_0 <= _GEN_497;
    end
    if (reset) begin
      vArrayWire_54_0 <= 1'h0;
    end else begin
      vArrayWire_54_0 <= _GEN_488;
    end
    if (reset) begin
      vArrayWire_53_0 <= 1'h0;
    end else begin
      vArrayWire_53_0 <= _GEN_479;
    end
    if (reset) begin
      vArrayWire_52_0 <= 1'h0;
    end else begin
      vArrayWire_52_0 <= _GEN_470;
    end
    if (reset) begin
      vArrayWire_51_0 <= 1'h0;
    end else begin
      vArrayWire_51_0 <= _GEN_461;
    end
    if (reset) begin
      vArrayWire_50_0 <= 1'h0;
    end else begin
      vArrayWire_50_0 <= _GEN_452;
    end
    if (reset) begin
      vArrayWire_49_0 <= 1'h0;
    end else begin
      vArrayWire_49_0 <= _GEN_443;
    end
    if (reset) begin
      vArrayWire_48_0 <= 1'h0;
    end else begin
      vArrayWire_48_0 <= _GEN_434;
    end
    if (reset) begin
      vArrayWire_47_0 <= 1'h0;
    end else begin
      vArrayWire_47_0 <= _GEN_425;
    end
    if (reset) begin
      vArrayWire_46_0 <= 1'h0;
    end else begin
      vArrayWire_46_0 <= _GEN_416;
    end
    if (reset) begin
      vArrayWire_45_0 <= 1'h0;
    end else begin
      vArrayWire_45_0 <= _GEN_407;
    end
    if (reset) begin
      vArrayWire_44_0 <= 1'h0;
    end else begin
      vArrayWire_44_0 <= _GEN_398;
    end
    if (reset) begin
      vArrayWire_43_0 <= 1'h0;
    end else begin
      vArrayWire_43_0 <= _GEN_389;
    end
    if (reset) begin
      vArrayWire_42_0 <= 1'h0;
    end else begin
      vArrayWire_42_0 <= _GEN_380;
    end
    if (reset) begin
      vArrayWire_41_0 <= 1'h0;
    end else begin
      vArrayWire_41_0 <= _GEN_371;
    end
    if (reset) begin
      vArrayWire_40_0 <= 1'h0;
    end else begin
      vArrayWire_40_0 <= _GEN_362;
    end
    if (reset) begin
      vArrayWire_39_0 <= 1'h0;
    end else begin
      vArrayWire_39_0 <= _GEN_353;
    end
    if (reset) begin
      vArrayWire_38_0 <= 1'h0;
    end else begin
      vArrayWire_38_0 <= _GEN_344;
    end
    if (reset) begin
      vArrayWire_37_0 <= 1'h0;
    end else begin
      vArrayWire_37_0 <= _GEN_335;
    end
    if (reset) begin
      vArrayWire_36_0 <= 1'h0;
    end else begin
      vArrayWire_36_0 <= _GEN_326;
    end
    if (reset) begin
      vArrayWire_35_0 <= 1'h0;
    end else begin
      vArrayWire_35_0 <= _GEN_317;
    end
    if (reset) begin
      vArrayWire_34_0 <= 1'h0;
    end else begin
      vArrayWire_34_0 <= _GEN_308;
    end
    if (reset) begin
      vArrayWire_33_0 <= 1'h0;
    end else begin
      vArrayWire_33_0 <= _GEN_299;
    end
    if (reset) begin
      vArrayWire_32_0 <= 1'h0;
    end else begin
      vArrayWire_32_0 <= _GEN_290;
    end
    if (reset) begin
      vArrayWire_31_0 <= 1'h0;
    end else begin
      vArrayWire_31_0 <= _GEN_281;
    end
    if (reset) begin
      vArrayWire_30_0 <= 1'h0;
    end else begin
      vArrayWire_30_0 <= _GEN_272;
    end
    if (reset) begin
      vArrayWire_29_0 <= 1'h0;
    end else begin
      vArrayWire_29_0 <= _GEN_263;
    end
    if (reset) begin
      vArrayWire_28_0 <= 1'h0;
    end else begin
      vArrayWire_28_0 <= _GEN_254;
    end
    if (reset) begin
      vArrayWire_27_0 <= 1'h0;
    end else begin
      vArrayWire_27_0 <= _GEN_245;
    end
    if (reset) begin
      vArrayWire_26_0 <= 1'h0;
    end else begin
      vArrayWire_26_0 <= _GEN_236;
    end
    if (reset) begin
      vArrayWire_25_0 <= 1'h0;
    end else begin
      vArrayWire_25_0 <= _GEN_227;
    end
    if (reset) begin
      vArrayWire_24_0 <= 1'h0;
    end else begin
      vArrayWire_24_0 <= _GEN_218;
    end
    if (reset) begin
      vArrayWire_23_0 <= 1'h0;
    end else begin
      vArrayWire_23_0 <= _GEN_209;
    end
    if (reset) begin
      vArrayWire_22_0 <= 1'h0;
    end else begin
      vArrayWire_22_0 <= _GEN_200;
    end
    if (reset) begin
      vArrayWire_21_0 <= 1'h0;
    end else begin
      vArrayWire_21_0 <= _GEN_191;
    end
    if (reset) begin
      vArrayWire_20_0 <= 1'h0;
    end else begin
      vArrayWire_20_0 <= _GEN_182;
    end
    if (reset) begin
      vArrayWire_19_0 <= 1'h0;
    end else begin
      vArrayWire_19_0 <= _GEN_173;
    end
    if (reset) begin
      vArrayWire_18_0 <= 1'h0;
    end else begin
      vArrayWire_18_0 <= _GEN_164;
    end
    if (reset) begin
      vArrayWire_17_0 <= 1'h0;
    end else begin
      vArrayWire_17_0 <= _GEN_155;
    end
    if (reset) begin
      vArrayWire_16_0 <= 1'h0;
    end else begin
      vArrayWire_16_0 <= _GEN_146;
    end
    if (reset) begin
      vArrayWire_15_0 <= 1'h0;
    end else begin
      vArrayWire_15_0 <= _GEN_137;
    end
    if (reset) begin
      vArrayWire_14_0 <= 1'h0;
    end else begin
      vArrayWire_14_0 <= _GEN_128;
    end
    if (reset) begin
      vArrayWire_13_0 <= 1'h0;
    end else begin
      vArrayWire_13_0 <= _GEN_119;
    end
    if (reset) begin
      vArrayWire_12_0 <= 1'h0;
    end else begin
      vArrayWire_12_0 <= _GEN_110;
    end
    if (reset) begin
      vArrayWire_11_0 <= 1'h0;
    end else begin
      vArrayWire_11_0 <= _GEN_101;
    end
    if (reset) begin
      vArrayWire_10_0 <= 1'h0;
    end else begin
      vArrayWire_10_0 <= _GEN_92;
    end
    if (reset) begin
      vArrayWire_9_0 <= 1'h0;
    end else begin
      vArrayWire_9_0 <= _GEN_83;
    end
    if (reset) begin
      vArrayWire_8_0 <= 1'h0;
    end else begin
      vArrayWire_8_0 <= _GEN_74;
    end
    if (reset) begin
      vArrayWire_7_0 <= 1'h0;
    end else begin
      vArrayWire_7_0 <= _GEN_65;
    end
    if (reset) begin
      vArrayWire_6_0 <= 1'h0;
    end else begin
      vArrayWire_6_0 <= _GEN_56;
    end
    if (reset) begin
      vArrayWire_5_0 <= 1'h0;
    end else begin
      vArrayWire_5_0 <= _GEN_47;
    end
    if (reset) begin
      vArrayWire_4_0 <= 1'h0;
    end else begin
      vArrayWire_4_0 <= _GEN_38;
    end
    if (reset) begin
      vArrayWire_3_0 <= 1'h0;
    end else begin
      vArrayWire_3_0 <= _GEN_29;
    end
    if (reset) begin
      vArrayWire_2_0 <= 1'h0;
    end else begin
      vArrayWire_2_0 <= _GEN_20;
    end
    if (reset) begin
      vArrayWire_1_0 <= 1'h0;
    end else begin
      vArrayWire_1_0 <= _GEN_11;
    end
    if (reset) begin
      vArrayWire_0_0 <= 1'h0;
    end else begin
      vArrayWire_0_0 <= _GEN_2;
    end
    if (reset) begin
      tagArrayWire_63_0 <= 22'h0;
    end else if (_T_3755) begin
      tagArrayWire_63_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_0 <= 22'h0;
    end else if (_T_3702) begin
      tagArrayWire_62_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_0 <= 22'h0;
    end else if (_T_3649) begin
      tagArrayWire_61_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_0 <= 22'h0;
    end else if (_T_3596) begin
      tagArrayWire_60_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_0 <= 22'h0;
    end else if (_T_3543) begin
      tagArrayWire_59_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_0 <= 22'h0;
    end else if (_T_3490) begin
      tagArrayWire_58_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_0 <= 22'h0;
    end else if (_T_3437) begin
      tagArrayWire_57_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_0 <= 22'h0;
    end else if (_T_3384) begin
      tagArrayWire_56_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_0 <= 22'h0;
    end else if (_T_3331) begin
      tagArrayWire_55_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_0 <= 22'h0;
    end else if (_T_3278) begin
      tagArrayWire_54_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_0 <= 22'h0;
    end else if (_T_3225) begin
      tagArrayWire_53_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_0 <= 22'h0;
    end else if (_T_3172) begin
      tagArrayWire_52_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_0 <= 22'h0;
    end else if (_T_3119) begin
      tagArrayWire_51_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_0 <= 22'h0;
    end else if (_T_3066) begin
      tagArrayWire_50_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_0 <= 22'h0;
    end else if (_T_3013) begin
      tagArrayWire_49_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_0 <= 22'h0;
    end else if (_T_2960) begin
      tagArrayWire_48_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_0 <= 22'h0;
    end else if (_T_2907) begin
      tagArrayWire_47_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_0 <= 22'h0;
    end else if (_T_2854) begin
      tagArrayWire_46_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_0 <= 22'h0;
    end else if (_T_2801) begin
      tagArrayWire_45_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_0 <= 22'h0;
    end else if (_T_2748) begin
      tagArrayWire_44_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_0 <= 22'h0;
    end else if (_T_2695) begin
      tagArrayWire_43_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_0 <= 22'h0;
    end else if (_T_2642) begin
      tagArrayWire_42_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_0 <= 22'h0;
    end else if (_T_2589) begin
      tagArrayWire_41_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_0 <= 22'h0;
    end else if (_T_2536) begin
      tagArrayWire_40_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_0 <= 22'h0;
    end else if (_T_2483) begin
      tagArrayWire_39_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_0 <= 22'h0;
    end else if (_T_2430) begin
      tagArrayWire_38_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_0 <= 22'h0;
    end else if (_T_2377) begin
      tagArrayWire_37_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_0 <= 22'h0;
    end else if (_T_2324) begin
      tagArrayWire_36_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_0 <= 22'h0;
    end else if (_T_2271) begin
      tagArrayWire_35_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_0 <= 22'h0;
    end else if (_T_2218) begin
      tagArrayWire_34_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_0 <= 22'h0;
    end else if (_T_2165) begin
      tagArrayWire_33_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_0 <= 22'h0;
    end else if (_T_2112) begin
      tagArrayWire_32_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_0 <= 22'h0;
    end else if (_T_2059) begin
      tagArrayWire_31_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_0 <= 22'h0;
    end else if (_T_2006) begin
      tagArrayWire_30_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_0 <= 22'h0;
    end else if (_T_1953) begin
      tagArrayWire_29_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_0 <= 22'h0;
    end else if (_T_1900) begin
      tagArrayWire_28_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_0 <= 22'h0;
    end else if (_T_1847) begin
      tagArrayWire_27_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_0 <= 22'h0;
    end else if (_T_1794) begin
      tagArrayWire_26_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_0 <= 22'h0;
    end else if (_T_1741) begin
      tagArrayWire_25_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_0 <= 22'h0;
    end else if (_T_1688) begin
      tagArrayWire_24_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_0 <= 22'h0;
    end else if (_T_1635) begin
      tagArrayWire_23_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_0 <= 22'h0;
    end else if (_T_1582) begin
      tagArrayWire_22_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_0 <= 22'h0;
    end else if (_T_1529) begin
      tagArrayWire_21_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_0 <= 22'h0;
    end else if (_T_1476) begin
      tagArrayWire_20_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_0 <= 22'h0;
    end else if (_T_1423) begin
      tagArrayWire_19_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_0 <= 22'h0;
    end else if (_T_1370) begin
      tagArrayWire_18_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_0 <= 22'h0;
    end else if (_T_1317) begin
      tagArrayWire_17_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_0 <= 22'h0;
    end else if (_T_1264) begin
      tagArrayWire_16_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_0 <= 22'h0;
    end else if (_T_1211) begin
      tagArrayWire_15_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_0 <= 22'h0;
    end else if (_T_1158) begin
      tagArrayWire_14_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_0 <= 22'h0;
    end else if (_T_1105) begin
      tagArrayWire_13_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_0 <= 22'h0;
    end else if (_T_1052) begin
      tagArrayWire_12_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_0 <= 22'h0;
    end else if (_T_999) begin
      tagArrayWire_11_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_0 <= 22'h0;
    end else if (_T_946) begin
      tagArrayWire_10_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_0 <= 22'h0;
    end else if (_T_893) begin
      tagArrayWire_9_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_0 <= 22'h0;
    end else if (_T_840) begin
      tagArrayWire_8_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_0 <= 22'h0;
    end else if (_T_787) begin
      tagArrayWire_7_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_0 <= 22'h0;
    end else if (_T_734) begin
      tagArrayWire_6_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_0 <= 22'h0;
    end else if (_T_681) begin
      tagArrayWire_5_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_0 <= 22'h0;
    end else if (_T_628) begin
      tagArrayWire_4_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_0 <= 22'h0;
    end else if (_T_575) begin
      tagArrayWire_3_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_0 <= 22'h0;
    end else if (_T_522) begin
      tagArrayWire_2_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_0 <= 22'h0;
    end else if (_T_469) begin
      tagArrayWire_1_0 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_0 <= 22'h0;
    end else if (_T_416) begin
      tagArrayWire_0_0 <= tag;
    end
    if (reset) begin
      vArrayWire_63_1 <= 1'h0;
    end else begin
      vArrayWire_63_1 <= _GEN_571;
    end
    if (reset) begin
      vArrayWire_62_1 <= 1'h0;
    end else begin
      vArrayWire_62_1 <= _GEN_562;
    end
    if (reset) begin
      vArrayWire_61_1 <= 1'h0;
    end else begin
      vArrayWire_61_1 <= _GEN_553;
    end
    if (reset) begin
      vArrayWire_60_1 <= 1'h0;
    end else begin
      vArrayWire_60_1 <= _GEN_544;
    end
    if (reset) begin
      vArrayWire_59_1 <= 1'h0;
    end else begin
      vArrayWire_59_1 <= _GEN_535;
    end
    if (reset) begin
      vArrayWire_58_1 <= 1'h0;
    end else begin
      vArrayWire_58_1 <= _GEN_526;
    end
    if (reset) begin
      vArrayWire_57_1 <= 1'h0;
    end else begin
      vArrayWire_57_1 <= _GEN_517;
    end
    if (reset) begin
      vArrayWire_56_1 <= 1'h0;
    end else begin
      vArrayWire_56_1 <= _GEN_508;
    end
    if (reset) begin
      vArrayWire_55_1 <= 1'h0;
    end else begin
      vArrayWire_55_1 <= _GEN_499;
    end
    if (reset) begin
      vArrayWire_54_1 <= 1'h0;
    end else begin
      vArrayWire_54_1 <= _GEN_490;
    end
    if (reset) begin
      vArrayWire_53_1 <= 1'h0;
    end else begin
      vArrayWire_53_1 <= _GEN_481;
    end
    if (reset) begin
      vArrayWire_52_1 <= 1'h0;
    end else begin
      vArrayWire_52_1 <= _GEN_472;
    end
    if (reset) begin
      vArrayWire_51_1 <= 1'h0;
    end else begin
      vArrayWire_51_1 <= _GEN_463;
    end
    if (reset) begin
      vArrayWire_50_1 <= 1'h0;
    end else begin
      vArrayWire_50_1 <= _GEN_454;
    end
    if (reset) begin
      vArrayWire_49_1 <= 1'h0;
    end else begin
      vArrayWire_49_1 <= _GEN_445;
    end
    if (reset) begin
      vArrayWire_48_1 <= 1'h0;
    end else begin
      vArrayWire_48_1 <= _GEN_436;
    end
    if (reset) begin
      vArrayWire_47_1 <= 1'h0;
    end else begin
      vArrayWire_47_1 <= _GEN_427;
    end
    if (reset) begin
      vArrayWire_46_1 <= 1'h0;
    end else begin
      vArrayWire_46_1 <= _GEN_418;
    end
    if (reset) begin
      vArrayWire_45_1 <= 1'h0;
    end else begin
      vArrayWire_45_1 <= _GEN_409;
    end
    if (reset) begin
      vArrayWire_44_1 <= 1'h0;
    end else begin
      vArrayWire_44_1 <= _GEN_400;
    end
    if (reset) begin
      vArrayWire_43_1 <= 1'h0;
    end else begin
      vArrayWire_43_1 <= _GEN_391;
    end
    if (reset) begin
      vArrayWire_42_1 <= 1'h0;
    end else begin
      vArrayWire_42_1 <= _GEN_382;
    end
    if (reset) begin
      vArrayWire_41_1 <= 1'h0;
    end else begin
      vArrayWire_41_1 <= _GEN_373;
    end
    if (reset) begin
      vArrayWire_40_1 <= 1'h0;
    end else begin
      vArrayWire_40_1 <= _GEN_364;
    end
    if (reset) begin
      vArrayWire_39_1 <= 1'h0;
    end else begin
      vArrayWire_39_1 <= _GEN_355;
    end
    if (reset) begin
      vArrayWire_38_1 <= 1'h0;
    end else begin
      vArrayWire_38_1 <= _GEN_346;
    end
    if (reset) begin
      vArrayWire_37_1 <= 1'h0;
    end else begin
      vArrayWire_37_1 <= _GEN_337;
    end
    if (reset) begin
      vArrayWire_36_1 <= 1'h0;
    end else begin
      vArrayWire_36_1 <= _GEN_328;
    end
    if (reset) begin
      vArrayWire_35_1 <= 1'h0;
    end else begin
      vArrayWire_35_1 <= _GEN_319;
    end
    if (reset) begin
      vArrayWire_34_1 <= 1'h0;
    end else begin
      vArrayWire_34_1 <= _GEN_310;
    end
    if (reset) begin
      vArrayWire_33_1 <= 1'h0;
    end else begin
      vArrayWire_33_1 <= _GEN_301;
    end
    if (reset) begin
      vArrayWire_32_1 <= 1'h0;
    end else begin
      vArrayWire_32_1 <= _GEN_292;
    end
    if (reset) begin
      vArrayWire_31_1 <= 1'h0;
    end else begin
      vArrayWire_31_1 <= _GEN_283;
    end
    if (reset) begin
      vArrayWire_30_1 <= 1'h0;
    end else begin
      vArrayWire_30_1 <= _GEN_274;
    end
    if (reset) begin
      vArrayWire_29_1 <= 1'h0;
    end else begin
      vArrayWire_29_1 <= _GEN_265;
    end
    if (reset) begin
      vArrayWire_28_1 <= 1'h0;
    end else begin
      vArrayWire_28_1 <= _GEN_256;
    end
    if (reset) begin
      vArrayWire_27_1 <= 1'h0;
    end else begin
      vArrayWire_27_1 <= _GEN_247;
    end
    if (reset) begin
      vArrayWire_26_1 <= 1'h0;
    end else begin
      vArrayWire_26_1 <= _GEN_238;
    end
    if (reset) begin
      vArrayWire_25_1 <= 1'h0;
    end else begin
      vArrayWire_25_1 <= _GEN_229;
    end
    if (reset) begin
      vArrayWire_24_1 <= 1'h0;
    end else begin
      vArrayWire_24_1 <= _GEN_220;
    end
    if (reset) begin
      vArrayWire_23_1 <= 1'h0;
    end else begin
      vArrayWire_23_1 <= _GEN_211;
    end
    if (reset) begin
      vArrayWire_22_1 <= 1'h0;
    end else begin
      vArrayWire_22_1 <= _GEN_202;
    end
    if (reset) begin
      vArrayWire_21_1 <= 1'h0;
    end else begin
      vArrayWire_21_1 <= _GEN_193;
    end
    if (reset) begin
      vArrayWire_20_1 <= 1'h0;
    end else begin
      vArrayWire_20_1 <= _GEN_184;
    end
    if (reset) begin
      vArrayWire_19_1 <= 1'h0;
    end else begin
      vArrayWire_19_1 <= _GEN_175;
    end
    if (reset) begin
      vArrayWire_18_1 <= 1'h0;
    end else begin
      vArrayWire_18_1 <= _GEN_166;
    end
    if (reset) begin
      vArrayWire_17_1 <= 1'h0;
    end else begin
      vArrayWire_17_1 <= _GEN_157;
    end
    if (reset) begin
      vArrayWire_16_1 <= 1'h0;
    end else begin
      vArrayWire_16_1 <= _GEN_148;
    end
    if (reset) begin
      vArrayWire_15_1 <= 1'h0;
    end else begin
      vArrayWire_15_1 <= _GEN_139;
    end
    if (reset) begin
      vArrayWire_14_1 <= 1'h0;
    end else begin
      vArrayWire_14_1 <= _GEN_130;
    end
    if (reset) begin
      vArrayWire_13_1 <= 1'h0;
    end else begin
      vArrayWire_13_1 <= _GEN_121;
    end
    if (reset) begin
      vArrayWire_12_1 <= 1'h0;
    end else begin
      vArrayWire_12_1 <= _GEN_112;
    end
    if (reset) begin
      vArrayWire_11_1 <= 1'h0;
    end else begin
      vArrayWire_11_1 <= _GEN_103;
    end
    if (reset) begin
      vArrayWire_10_1 <= 1'h0;
    end else begin
      vArrayWire_10_1 <= _GEN_94;
    end
    if (reset) begin
      vArrayWire_9_1 <= 1'h0;
    end else begin
      vArrayWire_9_1 <= _GEN_85;
    end
    if (reset) begin
      vArrayWire_8_1 <= 1'h0;
    end else begin
      vArrayWire_8_1 <= _GEN_76;
    end
    if (reset) begin
      vArrayWire_7_1 <= 1'h0;
    end else begin
      vArrayWire_7_1 <= _GEN_67;
    end
    if (reset) begin
      vArrayWire_6_1 <= 1'h0;
    end else begin
      vArrayWire_6_1 <= _GEN_58;
    end
    if (reset) begin
      vArrayWire_5_1 <= 1'h0;
    end else begin
      vArrayWire_5_1 <= _GEN_49;
    end
    if (reset) begin
      vArrayWire_4_1 <= 1'h0;
    end else begin
      vArrayWire_4_1 <= _GEN_40;
    end
    if (reset) begin
      vArrayWire_3_1 <= 1'h0;
    end else begin
      vArrayWire_3_1 <= _GEN_31;
    end
    if (reset) begin
      vArrayWire_2_1 <= 1'h0;
    end else begin
      vArrayWire_2_1 <= _GEN_22;
    end
    if (reset) begin
      vArrayWire_1_1 <= 1'h0;
    end else begin
      vArrayWire_1_1 <= _GEN_13;
    end
    if (reset) begin
      vArrayWire_0_1 <= 1'h0;
    end else begin
      vArrayWire_0_1 <= _GEN_4;
    end
    if (reset) begin
      tagArrayWire_63_1 <= 22'h0;
    end else if (_T_3767) begin
      tagArrayWire_63_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_1 <= 22'h0;
    end else if (_T_3714) begin
      tagArrayWire_62_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_1 <= 22'h0;
    end else if (_T_3661) begin
      tagArrayWire_61_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_1 <= 22'h0;
    end else if (_T_3608) begin
      tagArrayWire_60_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_1 <= 22'h0;
    end else if (_T_3555) begin
      tagArrayWire_59_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_1 <= 22'h0;
    end else if (_T_3502) begin
      tagArrayWire_58_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_1 <= 22'h0;
    end else if (_T_3449) begin
      tagArrayWire_57_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_1 <= 22'h0;
    end else if (_T_3396) begin
      tagArrayWire_56_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_1 <= 22'h0;
    end else if (_T_3343) begin
      tagArrayWire_55_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_1 <= 22'h0;
    end else if (_T_3290) begin
      tagArrayWire_54_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_1 <= 22'h0;
    end else if (_T_3237) begin
      tagArrayWire_53_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_1 <= 22'h0;
    end else if (_T_3184) begin
      tagArrayWire_52_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_1 <= 22'h0;
    end else if (_T_3131) begin
      tagArrayWire_51_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_1 <= 22'h0;
    end else if (_T_3078) begin
      tagArrayWire_50_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_1 <= 22'h0;
    end else if (_T_3025) begin
      tagArrayWire_49_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_1 <= 22'h0;
    end else if (_T_2972) begin
      tagArrayWire_48_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_1 <= 22'h0;
    end else if (_T_2919) begin
      tagArrayWire_47_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_1 <= 22'h0;
    end else if (_T_2866) begin
      tagArrayWire_46_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_1 <= 22'h0;
    end else if (_T_2813) begin
      tagArrayWire_45_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_1 <= 22'h0;
    end else if (_T_2760) begin
      tagArrayWire_44_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_1 <= 22'h0;
    end else if (_T_2707) begin
      tagArrayWire_43_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_1 <= 22'h0;
    end else if (_T_2654) begin
      tagArrayWire_42_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_1 <= 22'h0;
    end else if (_T_2601) begin
      tagArrayWire_41_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_1 <= 22'h0;
    end else if (_T_2548) begin
      tagArrayWire_40_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_1 <= 22'h0;
    end else if (_T_2495) begin
      tagArrayWire_39_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_1 <= 22'h0;
    end else if (_T_2442) begin
      tagArrayWire_38_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_1 <= 22'h0;
    end else if (_T_2389) begin
      tagArrayWire_37_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_1 <= 22'h0;
    end else if (_T_2336) begin
      tagArrayWire_36_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_1 <= 22'h0;
    end else if (_T_2283) begin
      tagArrayWire_35_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_1 <= 22'h0;
    end else if (_T_2230) begin
      tagArrayWire_34_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_1 <= 22'h0;
    end else if (_T_2177) begin
      tagArrayWire_33_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_1 <= 22'h0;
    end else if (_T_2124) begin
      tagArrayWire_32_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_1 <= 22'h0;
    end else if (_T_2071) begin
      tagArrayWire_31_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_1 <= 22'h0;
    end else if (_T_2018) begin
      tagArrayWire_30_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_1 <= 22'h0;
    end else if (_T_1965) begin
      tagArrayWire_29_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_1 <= 22'h0;
    end else if (_T_1912) begin
      tagArrayWire_28_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_1 <= 22'h0;
    end else if (_T_1859) begin
      tagArrayWire_27_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_1 <= 22'h0;
    end else if (_T_1806) begin
      tagArrayWire_26_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_1 <= 22'h0;
    end else if (_T_1753) begin
      tagArrayWire_25_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_1 <= 22'h0;
    end else if (_T_1700) begin
      tagArrayWire_24_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_1 <= 22'h0;
    end else if (_T_1647) begin
      tagArrayWire_23_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_1 <= 22'h0;
    end else if (_T_1594) begin
      tagArrayWire_22_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_1 <= 22'h0;
    end else if (_T_1541) begin
      tagArrayWire_21_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_1 <= 22'h0;
    end else if (_T_1488) begin
      tagArrayWire_20_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_1 <= 22'h0;
    end else if (_T_1435) begin
      tagArrayWire_19_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_1 <= 22'h0;
    end else if (_T_1382) begin
      tagArrayWire_18_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_1 <= 22'h0;
    end else if (_T_1329) begin
      tagArrayWire_17_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_1 <= 22'h0;
    end else if (_T_1276) begin
      tagArrayWire_16_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_1 <= 22'h0;
    end else if (_T_1223) begin
      tagArrayWire_15_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_1 <= 22'h0;
    end else if (_T_1170) begin
      tagArrayWire_14_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_1 <= 22'h0;
    end else if (_T_1117) begin
      tagArrayWire_13_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_1 <= 22'h0;
    end else if (_T_1064) begin
      tagArrayWire_12_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_1 <= 22'h0;
    end else if (_T_1011) begin
      tagArrayWire_11_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_1 <= 22'h0;
    end else if (_T_958) begin
      tagArrayWire_10_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_1 <= 22'h0;
    end else if (_T_905) begin
      tagArrayWire_9_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_1 <= 22'h0;
    end else if (_T_852) begin
      tagArrayWire_8_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_1 <= 22'h0;
    end else if (_T_799) begin
      tagArrayWire_7_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_1 <= 22'h0;
    end else if (_T_746) begin
      tagArrayWire_6_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_1 <= 22'h0;
    end else if (_T_693) begin
      tagArrayWire_5_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_1 <= 22'h0;
    end else if (_T_640) begin
      tagArrayWire_4_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_1 <= 22'h0;
    end else if (_T_587) begin
      tagArrayWire_3_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_1 <= 22'h0;
    end else if (_T_534) begin
      tagArrayWire_2_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_1 <= 22'h0;
    end else if (_T_481) begin
      tagArrayWire_1_1 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_1 <= 22'h0;
    end else if (_T_428) begin
      tagArrayWire_0_1 <= tag;
    end
    if (reset) begin
      vArrayWire_63_2 <= 1'h0;
    end else begin
      vArrayWire_63_2 <= _GEN_573;
    end
    if (reset) begin
      vArrayWire_62_2 <= 1'h0;
    end else begin
      vArrayWire_62_2 <= _GEN_564;
    end
    if (reset) begin
      vArrayWire_61_2 <= 1'h0;
    end else begin
      vArrayWire_61_2 <= _GEN_555;
    end
    if (reset) begin
      vArrayWire_60_2 <= 1'h0;
    end else begin
      vArrayWire_60_2 <= _GEN_546;
    end
    if (reset) begin
      vArrayWire_59_2 <= 1'h0;
    end else begin
      vArrayWire_59_2 <= _GEN_537;
    end
    if (reset) begin
      vArrayWire_58_2 <= 1'h0;
    end else begin
      vArrayWire_58_2 <= _GEN_528;
    end
    if (reset) begin
      vArrayWire_57_2 <= 1'h0;
    end else begin
      vArrayWire_57_2 <= _GEN_519;
    end
    if (reset) begin
      vArrayWire_56_2 <= 1'h0;
    end else begin
      vArrayWire_56_2 <= _GEN_510;
    end
    if (reset) begin
      vArrayWire_55_2 <= 1'h0;
    end else begin
      vArrayWire_55_2 <= _GEN_501;
    end
    if (reset) begin
      vArrayWire_54_2 <= 1'h0;
    end else begin
      vArrayWire_54_2 <= _GEN_492;
    end
    if (reset) begin
      vArrayWire_53_2 <= 1'h0;
    end else begin
      vArrayWire_53_2 <= _GEN_483;
    end
    if (reset) begin
      vArrayWire_52_2 <= 1'h0;
    end else begin
      vArrayWire_52_2 <= _GEN_474;
    end
    if (reset) begin
      vArrayWire_51_2 <= 1'h0;
    end else begin
      vArrayWire_51_2 <= _GEN_465;
    end
    if (reset) begin
      vArrayWire_50_2 <= 1'h0;
    end else begin
      vArrayWire_50_2 <= _GEN_456;
    end
    if (reset) begin
      vArrayWire_49_2 <= 1'h0;
    end else begin
      vArrayWire_49_2 <= _GEN_447;
    end
    if (reset) begin
      vArrayWire_48_2 <= 1'h0;
    end else begin
      vArrayWire_48_2 <= _GEN_438;
    end
    if (reset) begin
      vArrayWire_47_2 <= 1'h0;
    end else begin
      vArrayWire_47_2 <= _GEN_429;
    end
    if (reset) begin
      vArrayWire_46_2 <= 1'h0;
    end else begin
      vArrayWire_46_2 <= _GEN_420;
    end
    if (reset) begin
      vArrayWire_45_2 <= 1'h0;
    end else begin
      vArrayWire_45_2 <= _GEN_411;
    end
    if (reset) begin
      vArrayWire_44_2 <= 1'h0;
    end else begin
      vArrayWire_44_2 <= _GEN_402;
    end
    if (reset) begin
      vArrayWire_43_2 <= 1'h0;
    end else begin
      vArrayWire_43_2 <= _GEN_393;
    end
    if (reset) begin
      vArrayWire_42_2 <= 1'h0;
    end else begin
      vArrayWire_42_2 <= _GEN_384;
    end
    if (reset) begin
      vArrayWire_41_2 <= 1'h0;
    end else begin
      vArrayWire_41_2 <= _GEN_375;
    end
    if (reset) begin
      vArrayWire_40_2 <= 1'h0;
    end else begin
      vArrayWire_40_2 <= _GEN_366;
    end
    if (reset) begin
      vArrayWire_39_2 <= 1'h0;
    end else begin
      vArrayWire_39_2 <= _GEN_357;
    end
    if (reset) begin
      vArrayWire_38_2 <= 1'h0;
    end else begin
      vArrayWire_38_2 <= _GEN_348;
    end
    if (reset) begin
      vArrayWire_37_2 <= 1'h0;
    end else begin
      vArrayWire_37_2 <= _GEN_339;
    end
    if (reset) begin
      vArrayWire_36_2 <= 1'h0;
    end else begin
      vArrayWire_36_2 <= _GEN_330;
    end
    if (reset) begin
      vArrayWire_35_2 <= 1'h0;
    end else begin
      vArrayWire_35_2 <= _GEN_321;
    end
    if (reset) begin
      vArrayWire_34_2 <= 1'h0;
    end else begin
      vArrayWire_34_2 <= _GEN_312;
    end
    if (reset) begin
      vArrayWire_33_2 <= 1'h0;
    end else begin
      vArrayWire_33_2 <= _GEN_303;
    end
    if (reset) begin
      vArrayWire_32_2 <= 1'h0;
    end else begin
      vArrayWire_32_2 <= _GEN_294;
    end
    if (reset) begin
      vArrayWire_31_2 <= 1'h0;
    end else begin
      vArrayWire_31_2 <= _GEN_285;
    end
    if (reset) begin
      vArrayWire_30_2 <= 1'h0;
    end else begin
      vArrayWire_30_2 <= _GEN_276;
    end
    if (reset) begin
      vArrayWire_29_2 <= 1'h0;
    end else begin
      vArrayWire_29_2 <= _GEN_267;
    end
    if (reset) begin
      vArrayWire_28_2 <= 1'h0;
    end else begin
      vArrayWire_28_2 <= _GEN_258;
    end
    if (reset) begin
      vArrayWire_27_2 <= 1'h0;
    end else begin
      vArrayWire_27_2 <= _GEN_249;
    end
    if (reset) begin
      vArrayWire_26_2 <= 1'h0;
    end else begin
      vArrayWire_26_2 <= _GEN_240;
    end
    if (reset) begin
      vArrayWire_25_2 <= 1'h0;
    end else begin
      vArrayWire_25_2 <= _GEN_231;
    end
    if (reset) begin
      vArrayWire_24_2 <= 1'h0;
    end else begin
      vArrayWire_24_2 <= _GEN_222;
    end
    if (reset) begin
      vArrayWire_23_2 <= 1'h0;
    end else begin
      vArrayWire_23_2 <= _GEN_213;
    end
    if (reset) begin
      vArrayWire_22_2 <= 1'h0;
    end else begin
      vArrayWire_22_2 <= _GEN_204;
    end
    if (reset) begin
      vArrayWire_21_2 <= 1'h0;
    end else begin
      vArrayWire_21_2 <= _GEN_195;
    end
    if (reset) begin
      vArrayWire_20_2 <= 1'h0;
    end else begin
      vArrayWire_20_2 <= _GEN_186;
    end
    if (reset) begin
      vArrayWire_19_2 <= 1'h0;
    end else begin
      vArrayWire_19_2 <= _GEN_177;
    end
    if (reset) begin
      vArrayWire_18_2 <= 1'h0;
    end else begin
      vArrayWire_18_2 <= _GEN_168;
    end
    if (reset) begin
      vArrayWire_17_2 <= 1'h0;
    end else begin
      vArrayWire_17_2 <= _GEN_159;
    end
    if (reset) begin
      vArrayWire_16_2 <= 1'h0;
    end else begin
      vArrayWire_16_2 <= _GEN_150;
    end
    if (reset) begin
      vArrayWire_15_2 <= 1'h0;
    end else begin
      vArrayWire_15_2 <= _GEN_141;
    end
    if (reset) begin
      vArrayWire_14_2 <= 1'h0;
    end else begin
      vArrayWire_14_2 <= _GEN_132;
    end
    if (reset) begin
      vArrayWire_13_2 <= 1'h0;
    end else begin
      vArrayWire_13_2 <= _GEN_123;
    end
    if (reset) begin
      vArrayWire_12_2 <= 1'h0;
    end else begin
      vArrayWire_12_2 <= _GEN_114;
    end
    if (reset) begin
      vArrayWire_11_2 <= 1'h0;
    end else begin
      vArrayWire_11_2 <= _GEN_105;
    end
    if (reset) begin
      vArrayWire_10_2 <= 1'h0;
    end else begin
      vArrayWire_10_2 <= _GEN_96;
    end
    if (reset) begin
      vArrayWire_9_2 <= 1'h0;
    end else begin
      vArrayWire_9_2 <= _GEN_87;
    end
    if (reset) begin
      vArrayWire_8_2 <= 1'h0;
    end else begin
      vArrayWire_8_2 <= _GEN_78;
    end
    if (reset) begin
      vArrayWire_7_2 <= 1'h0;
    end else begin
      vArrayWire_7_2 <= _GEN_69;
    end
    if (reset) begin
      vArrayWire_6_2 <= 1'h0;
    end else begin
      vArrayWire_6_2 <= _GEN_60;
    end
    if (reset) begin
      vArrayWire_5_2 <= 1'h0;
    end else begin
      vArrayWire_5_2 <= _GEN_51;
    end
    if (reset) begin
      vArrayWire_4_2 <= 1'h0;
    end else begin
      vArrayWire_4_2 <= _GEN_42;
    end
    if (reset) begin
      vArrayWire_3_2 <= 1'h0;
    end else begin
      vArrayWire_3_2 <= _GEN_33;
    end
    if (reset) begin
      vArrayWire_2_2 <= 1'h0;
    end else begin
      vArrayWire_2_2 <= _GEN_24;
    end
    if (reset) begin
      vArrayWire_1_2 <= 1'h0;
    end else begin
      vArrayWire_1_2 <= _GEN_15;
    end
    if (reset) begin
      vArrayWire_0_2 <= 1'h0;
    end else begin
      vArrayWire_0_2 <= _GEN_6;
    end
    if (reset) begin
      tagArrayWire_63_2 <= 22'h0;
    end else if (_T_3779) begin
      tagArrayWire_63_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_2 <= 22'h0;
    end else if (_T_3726) begin
      tagArrayWire_62_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_2 <= 22'h0;
    end else if (_T_3673) begin
      tagArrayWire_61_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_2 <= 22'h0;
    end else if (_T_3620) begin
      tagArrayWire_60_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_2 <= 22'h0;
    end else if (_T_3567) begin
      tagArrayWire_59_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_2 <= 22'h0;
    end else if (_T_3514) begin
      tagArrayWire_58_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_2 <= 22'h0;
    end else if (_T_3461) begin
      tagArrayWire_57_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_2 <= 22'h0;
    end else if (_T_3408) begin
      tagArrayWire_56_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_2 <= 22'h0;
    end else if (_T_3355) begin
      tagArrayWire_55_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_2 <= 22'h0;
    end else if (_T_3302) begin
      tagArrayWire_54_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_2 <= 22'h0;
    end else if (_T_3249) begin
      tagArrayWire_53_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_2 <= 22'h0;
    end else if (_T_3196) begin
      tagArrayWire_52_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_2 <= 22'h0;
    end else if (_T_3143) begin
      tagArrayWire_51_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_2 <= 22'h0;
    end else if (_T_3090) begin
      tagArrayWire_50_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_2 <= 22'h0;
    end else if (_T_3037) begin
      tagArrayWire_49_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_2 <= 22'h0;
    end else if (_T_2984) begin
      tagArrayWire_48_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_2 <= 22'h0;
    end else if (_T_2931) begin
      tagArrayWire_47_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_2 <= 22'h0;
    end else if (_T_2878) begin
      tagArrayWire_46_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_2 <= 22'h0;
    end else if (_T_2825) begin
      tagArrayWire_45_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_2 <= 22'h0;
    end else if (_T_2772) begin
      tagArrayWire_44_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_2 <= 22'h0;
    end else if (_T_2719) begin
      tagArrayWire_43_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_2 <= 22'h0;
    end else if (_T_2666) begin
      tagArrayWire_42_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_2 <= 22'h0;
    end else if (_T_2613) begin
      tagArrayWire_41_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_2 <= 22'h0;
    end else if (_T_2560) begin
      tagArrayWire_40_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_2 <= 22'h0;
    end else if (_T_2507) begin
      tagArrayWire_39_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_2 <= 22'h0;
    end else if (_T_2454) begin
      tagArrayWire_38_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_2 <= 22'h0;
    end else if (_T_2401) begin
      tagArrayWire_37_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_2 <= 22'h0;
    end else if (_T_2348) begin
      tagArrayWire_36_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_2 <= 22'h0;
    end else if (_T_2295) begin
      tagArrayWire_35_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_2 <= 22'h0;
    end else if (_T_2242) begin
      tagArrayWire_34_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_2 <= 22'h0;
    end else if (_T_2189) begin
      tagArrayWire_33_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_2 <= 22'h0;
    end else if (_T_2136) begin
      tagArrayWire_32_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_2 <= 22'h0;
    end else if (_T_2083) begin
      tagArrayWire_31_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_2 <= 22'h0;
    end else if (_T_2030) begin
      tagArrayWire_30_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_2 <= 22'h0;
    end else if (_T_1977) begin
      tagArrayWire_29_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_2 <= 22'h0;
    end else if (_T_1924) begin
      tagArrayWire_28_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_2 <= 22'h0;
    end else if (_T_1871) begin
      tagArrayWire_27_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_2 <= 22'h0;
    end else if (_T_1818) begin
      tagArrayWire_26_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_2 <= 22'h0;
    end else if (_T_1765) begin
      tagArrayWire_25_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_2 <= 22'h0;
    end else if (_T_1712) begin
      tagArrayWire_24_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_2 <= 22'h0;
    end else if (_T_1659) begin
      tagArrayWire_23_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_2 <= 22'h0;
    end else if (_T_1606) begin
      tagArrayWire_22_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_2 <= 22'h0;
    end else if (_T_1553) begin
      tagArrayWire_21_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_2 <= 22'h0;
    end else if (_T_1500) begin
      tagArrayWire_20_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_2 <= 22'h0;
    end else if (_T_1447) begin
      tagArrayWire_19_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_2 <= 22'h0;
    end else if (_T_1394) begin
      tagArrayWire_18_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_2 <= 22'h0;
    end else if (_T_1341) begin
      tagArrayWire_17_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_2 <= 22'h0;
    end else if (_T_1288) begin
      tagArrayWire_16_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_2 <= 22'h0;
    end else if (_T_1235) begin
      tagArrayWire_15_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_2 <= 22'h0;
    end else if (_T_1182) begin
      tagArrayWire_14_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_2 <= 22'h0;
    end else if (_T_1129) begin
      tagArrayWire_13_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_2 <= 22'h0;
    end else if (_T_1076) begin
      tagArrayWire_12_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_2 <= 22'h0;
    end else if (_T_1023) begin
      tagArrayWire_11_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_2 <= 22'h0;
    end else if (_T_970) begin
      tagArrayWire_10_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_2 <= 22'h0;
    end else if (_T_917) begin
      tagArrayWire_9_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_2 <= 22'h0;
    end else if (_T_864) begin
      tagArrayWire_8_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_2 <= 22'h0;
    end else if (_T_811) begin
      tagArrayWire_7_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_2 <= 22'h0;
    end else if (_T_758) begin
      tagArrayWire_6_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_2 <= 22'h0;
    end else if (_T_705) begin
      tagArrayWire_5_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_2 <= 22'h0;
    end else if (_T_652) begin
      tagArrayWire_4_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_2 <= 22'h0;
    end else if (_T_599) begin
      tagArrayWire_3_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_2 <= 22'h0;
    end else if (_T_546) begin
      tagArrayWire_2_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_2 <= 22'h0;
    end else if (_T_493) begin
      tagArrayWire_1_2 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_2 <= 22'h0;
    end else if (_T_440) begin
      tagArrayWire_0_2 <= tag;
    end
    if (reset) begin
      vArrayWire_63_3 <= 1'h0;
    end else begin
      vArrayWire_63_3 <= _GEN_575;
    end
    if (reset) begin
      vArrayWire_62_3 <= 1'h0;
    end else begin
      vArrayWire_62_3 <= _GEN_566;
    end
    if (reset) begin
      vArrayWire_61_3 <= 1'h0;
    end else begin
      vArrayWire_61_3 <= _GEN_557;
    end
    if (reset) begin
      vArrayWire_60_3 <= 1'h0;
    end else begin
      vArrayWire_60_3 <= _GEN_548;
    end
    if (reset) begin
      vArrayWire_59_3 <= 1'h0;
    end else begin
      vArrayWire_59_3 <= _GEN_539;
    end
    if (reset) begin
      vArrayWire_58_3 <= 1'h0;
    end else begin
      vArrayWire_58_3 <= _GEN_530;
    end
    if (reset) begin
      vArrayWire_57_3 <= 1'h0;
    end else begin
      vArrayWire_57_3 <= _GEN_521;
    end
    if (reset) begin
      vArrayWire_56_3 <= 1'h0;
    end else begin
      vArrayWire_56_3 <= _GEN_512;
    end
    if (reset) begin
      vArrayWire_55_3 <= 1'h0;
    end else begin
      vArrayWire_55_3 <= _GEN_503;
    end
    if (reset) begin
      vArrayWire_54_3 <= 1'h0;
    end else begin
      vArrayWire_54_3 <= _GEN_494;
    end
    if (reset) begin
      vArrayWire_53_3 <= 1'h0;
    end else begin
      vArrayWire_53_3 <= _GEN_485;
    end
    if (reset) begin
      vArrayWire_52_3 <= 1'h0;
    end else begin
      vArrayWire_52_3 <= _GEN_476;
    end
    if (reset) begin
      vArrayWire_51_3 <= 1'h0;
    end else begin
      vArrayWire_51_3 <= _GEN_467;
    end
    if (reset) begin
      vArrayWire_50_3 <= 1'h0;
    end else begin
      vArrayWire_50_3 <= _GEN_458;
    end
    if (reset) begin
      vArrayWire_49_3 <= 1'h0;
    end else begin
      vArrayWire_49_3 <= _GEN_449;
    end
    if (reset) begin
      vArrayWire_48_3 <= 1'h0;
    end else begin
      vArrayWire_48_3 <= _GEN_440;
    end
    if (reset) begin
      vArrayWire_47_3 <= 1'h0;
    end else begin
      vArrayWire_47_3 <= _GEN_431;
    end
    if (reset) begin
      vArrayWire_46_3 <= 1'h0;
    end else begin
      vArrayWire_46_3 <= _GEN_422;
    end
    if (reset) begin
      vArrayWire_45_3 <= 1'h0;
    end else begin
      vArrayWire_45_3 <= _GEN_413;
    end
    if (reset) begin
      vArrayWire_44_3 <= 1'h0;
    end else begin
      vArrayWire_44_3 <= _GEN_404;
    end
    if (reset) begin
      vArrayWire_43_3 <= 1'h0;
    end else begin
      vArrayWire_43_3 <= _GEN_395;
    end
    if (reset) begin
      vArrayWire_42_3 <= 1'h0;
    end else begin
      vArrayWire_42_3 <= _GEN_386;
    end
    if (reset) begin
      vArrayWire_41_3 <= 1'h0;
    end else begin
      vArrayWire_41_3 <= _GEN_377;
    end
    if (reset) begin
      vArrayWire_40_3 <= 1'h0;
    end else begin
      vArrayWire_40_3 <= _GEN_368;
    end
    if (reset) begin
      vArrayWire_39_3 <= 1'h0;
    end else begin
      vArrayWire_39_3 <= _GEN_359;
    end
    if (reset) begin
      vArrayWire_38_3 <= 1'h0;
    end else begin
      vArrayWire_38_3 <= _GEN_350;
    end
    if (reset) begin
      vArrayWire_37_3 <= 1'h0;
    end else begin
      vArrayWire_37_3 <= _GEN_341;
    end
    if (reset) begin
      vArrayWire_36_3 <= 1'h0;
    end else begin
      vArrayWire_36_3 <= _GEN_332;
    end
    if (reset) begin
      vArrayWire_35_3 <= 1'h0;
    end else begin
      vArrayWire_35_3 <= _GEN_323;
    end
    if (reset) begin
      vArrayWire_34_3 <= 1'h0;
    end else begin
      vArrayWire_34_3 <= _GEN_314;
    end
    if (reset) begin
      vArrayWire_33_3 <= 1'h0;
    end else begin
      vArrayWire_33_3 <= _GEN_305;
    end
    if (reset) begin
      vArrayWire_32_3 <= 1'h0;
    end else begin
      vArrayWire_32_3 <= _GEN_296;
    end
    if (reset) begin
      vArrayWire_31_3 <= 1'h0;
    end else begin
      vArrayWire_31_3 <= _GEN_287;
    end
    if (reset) begin
      vArrayWire_30_3 <= 1'h0;
    end else begin
      vArrayWire_30_3 <= _GEN_278;
    end
    if (reset) begin
      vArrayWire_29_3 <= 1'h0;
    end else begin
      vArrayWire_29_3 <= _GEN_269;
    end
    if (reset) begin
      vArrayWire_28_3 <= 1'h0;
    end else begin
      vArrayWire_28_3 <= _GEN_260;
    end
    if (reset) begin
      vArrayWire_27_3 <= 1'h0;
    end else begin
      vArrayWire_27_3 <= _GEN_251;
    end
    if (reset) begin
      vArrayWire_26_3 <= 1'h0;
    end else begin
      vArrayWire_26_3 <= _GEN_242;
    end
    if (reset) begin
      vArrayWire_25_3 <= 1'h0;
    end else begin
      vArrayWire_25_3 <= _GEN_233;
    end
    if (reset) begin
      vArrayWire_24_3 <= 1'h0;
    end else begin
      vArrayWire_24_3 <= _GEN_224;
    end
    if (reset) begin
      vArrayWire_23_3 <= 1'h0;
    end else begin
      vArrayWire_23_3 <= _GEN_215;
    end
    if (reset) begin
      vArrayWire_22_3 <= 1'h0;
    end else begin
      vArrayWire_22_3 <= _GEN_206;
    end
    if (reset) begin
      vArrayWire_21_3 <= 1'h0;
    end else begin
      vArrayWire_21_3 <= _GEN_197;
    end
    if (reset) begin
      vArrayWire_20_3 <= 1'h0;
    end else begin
      vArrayWire_20_3 <= _GEN_188;
    end
    if (reset) begin
      vArrayWire_19_3 <= 1'h0;
    end else begin
      vArrayWire_19_3 <= _GEN_179;
    end
    if (reset) begin
      vArrayWire_18_3 <= 1'h0;
    end else begin
      vArrayWire_18_3 <= _GEN_170;
    end
    if (reset) begin
      vArrayWire_17_3 <= 1'h0;
    end else begin
      vArrayWire_17_3 <= _GEN_161;
    end
    if (reset) begin
      vArrayWire_16_3 <= 1'h0;
    end else begin
      vArrayWire_16_3 <= _GEN_152;
    end
    if (reset) begin
      vArrayWire_15_3 <= 1'h0;
    end else begin
      vArrayWire_15_3 <= _GEN_143;
    end
    if (reset) begin
      vArrayWire_14_3 <= 1'h0;
    end else begin
      vArrayWire_14_3 <= _GEN_134;
    end
    if (reset) begin
      vArrayWire_13_3 <= 1'h0;
    end else begin
      vArrayWire_13_3 <= _GEN_125;
    end
    if (reset) begin
      vArrayWire_12_3 <= 1'h0;
    end else begin
      vArrayWire_12_3 <= _GEN_116;
    end
    if (reset) begin
      vArrayWire_11_3 <= 1'h0;
    end else begin
      vArrayWire_11_3 <= _GEN_107;
    end
    if (reset) begin
      vArrayWire_10_3 <= 1'h0;
    end else begin
      vArrayWire_10_3 <= _GEN_98;
    end
    if (reset) begin
      vArrayWire_9_3 <= 1'h0;
    end else begin
      vArrayWire_9_3 <= _GEN_89;
    end
    if (reset) begin
      vArrayWire_8_3 <= 1'h0;
    end else begin
      vArrayWire_8_3 <= _GEN_80;
    end
    if (reset) begin
      vArrayWire_7_3 <= 1'h0;
    end else begin
      vArrayWire_7_3 <= _GEN_71;
    end
    if (reset) begin
      vArrayWire_6_3 <= 1'h0;
    end else begin
      vArrayWire_6_3 <= _GEN_62;
    end
    if (reset) begin
      vArrayWire_5_3 <= 1'h0;
    end else begin
      vArrayWire_5_3 <= _GEN_53;
    end
    if (reset) begin
      vArrayWire_4_3 <= 1'h0;
    end else begin
      vArrayWire_4_3 <= _GEN_44;
    end
    if (reset) begin
      vArrayWire_3_3 <= 1'h0;
    end else begin
      vArrayWire_3_3 <= _GEN_35;
    end
    if (reset) begin
      vArrayWire_2_3 <= 1'h0;
    end else begin
      vArrayWire_2_3 <= _GEN_26;
    end
    if (reset) begin
      vArrayWire_1_3 <= 1'h0;
    end else begin
      vArrayWire_1_3 <= _GEN_17;
    end
    if (reset) begin
      vArrayWire_0_3 <= 1'h0;
    end else begin
      vArrayWire_0_3 <= _GEN_8;
    end
    if (reset) begin
      tagArrayWire_63_3 <= 22'h0;
    end else if (_T_3791) begin
      tagArrayWire_63_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_62_3 <= 22'h0;
    end else if (_T_3738) begin
      tagArrayWire_62_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_61_3 <= 22'h0;
    end else if (_T_3685) begin
      tagArrayWire_61_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_60_3 <= 22'h0;
    end else if (_T_3632) begin
      tagArrayWire_60_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_59_3 <= 22'h0;
    end else if (_T_3579) begin
      tagArrayWire_59_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_58_3 <= 22'h0;
    end else if (_T_3526) begin
      tagArrayWire_58_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_57_3 <= 22'h0;
    end else if (_T_3473) begin
      tagArrayWire_57_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_56_3 <= 22'h0;
    end else if (_T_3420) begin
      tagArrayWire_56_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_55_3 <= 22'h0;
    end else if (_T_3367) begin
      tagArrayWire_55_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_54_3 <= 22'h0;
    end else if (_T_3314) begin
      tagArrayWire_54_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_53_3 <= 22'h0;
    end else if (_T_3261) begin
      tagArrayWire_53_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_52_3 <= 22'h0;
    end else if (_T_3208) begin
      tagArrayWire_52_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_51_3 <= 22'h0;
    end else if (_T_3155) begin
      tagArrayWire_51_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_50_3 <= 22'h0;
    end else if (_T_3102) begin
      tagArrayWire_50_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_49_3 <= 22'h0;
    end else if (_T_3049) begin
      tagArrayWire_49_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_48_3 <= 22'h0;
    end else if (_T_2996) begin
      tagArrayWire_48_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_47_3 <= 22'h0;
    end else if (_T_2943) begin
      tagArrayWire_47_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_46_3 <= 22'h0;
    end else if (_T_2890) begin
      tagArrayWire_46_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_45_3 <= 22'h0;
    end else if (_T_2837) begin
      tagArrayWire_45_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_44_3 <= 22'h0;
    end else if (_T_2784) begin
      tagArrayWire_44_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_43_3 <= 22'h0;
    end else if (_T_2731) begin
      tagArrayWire_43_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_42_3 <= 22'h0;
    end else if (_T_2678) begin
      tagArrayWire_42_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_41_3 <= 22'h0;
    end else if (_T_2625) begin
      tagArrayWire_41_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_40_3 <= 22'h0;
    end else if (_T_2572) begin
      tagArrayWire_40_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_39_3 <= 22'h0;
    end else if (_T_2519) begin
      tagArrayWire_39_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_38_3 <= 22'h0;
    end else if (_T_2466) begin
      tagArrayWire_38_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_37_3 <= 22'h0;
    end else if (_T_2413) begin
      tagArrayWire_37_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_36_3 <= 22'h0;
    end else if (_T_2360) begin
      tagArrayWire_36_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_35_3 <= 22'h0;
    end else if (_T_2307) begin
      tagArrayWire_35_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_34_3 <= 22'h0;
    end else if (_T_2254) begin
      tagArrayWire_34_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_33_3 <= 22'h0;
    end else if (_T_2201) begin
      tagArrayWire_33_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_32_3 <= 22'h0;
    end else if (_T_2148) begin
      tagArrayWire_32_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_31_3 <= 22'h0;
    end else if (_T_2095) begin
      tagArrayWire_31_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_30_3 <= 22'h0;
    end else if (_T_2042) begin
      tagArrayWire_30_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_29_3 <= 22'h0;
    end else if (_T_1989) begin
      tagArrayWire_29_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_28_3 <= 22'h0;
    end else if (_T_1936) begin
      tagArrayWire_28_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_27_3 <= 22'h0;
    end else if (_T_1883) begin
      tagArrayWire_27_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_26_3 <= 22'h0;
    end else if (_T_1830) begin
      tagArrayWire_26_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_25_3 <= 22'h0;
    end else if (_T_1777) begin
      tagArrayWire_25_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_24_3 <= 22'h0;
    end else if (_T_1724) begin
      tagArrayWire_24_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_23_3 <= 22'h0;
    end else if (_T_1671) begin
      tagArrayWire_23_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_22_3 <= 22'h0;
    end else if (_T_1618) begin
      tagArrayWire_22_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_21_3 <= 22'h0;
    end else if (_T_1565) begin
      tagArrayWire_21_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_20_3 <= 22'h0;
    end else if (_T_1512) begin
      tagArrayWire_20_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_19_3 <= 22'h0;
    end else if (_T_1459) begin
      tagArrayWire_19_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_18_3 <= 22'h0;
    end else if (_T_1406) begin
      tagArrayWire_18_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_17_3 <= 22'h0;
    end else if (_T_1353) begin
      tagArrayWire_17_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_16_3 <= 22'h0;
    end else if (_T_1300) begin
      tagArrayWire_16_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_15_3 <= 22'h0;
    end else if (_T_1247) begin
      tagArrayWire_15_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_14_3 <= 22'h0;
    end else if (_T_1194) begin
      tagArrayWire_14_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_13_3 <= 22'h0;
    end else if (_T_1141) begin
      tagArrayWire_13_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_12_3 <= 22'h0;
    end else if (_T_1088) begin
      tagArrayWire_12_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_11_3 <= 22'h0;
    end else if (_T_1035) begin
      tagArrayWire_11_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_10_3 <= 22'h0;
    end else if (_T_982) begin
      tagArrayWire_10_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_9_3 <= 22'h0;
    end else if (_T_929) begin
      tagArrayWire_9_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_8_3 <= 22'h0;
    end else if (_T_876) begin
      tagArrayWire_8_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_7_3 <= 22'h0;
    end else if (_T_823) begin
      tagArrayWire_7_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_6_3 <= 22'h0;
    end else if (_T_770) begin
      tagArrayWire_6_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_5_3 <= 22'h0;
    end else if (_T_717) begin
      tagArrayWire_5_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_4_3 <= 22'h0;
    end else if (_T_664) begin
      tagArrayWire_4_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_3_3 <= 22'h0;
    end else if (_T_611) begin
      tagArrayWire_3_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_2_3 <= 22'h0;
    end else if (_T_558) begin
      tagArrayWire_2_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_1_3 <= 22'h0;
    end else if (_T_505) begin
      tagArrayWire_1_3 <= tag;
    end
    if (reset) begin
      tagArrayWire_0_3 <= 22'h0;
    end else if (_T_452) begin
      tagArrayWire_0_3 <= tag;
    end
    if (reset) begin
      selArrayWire_1 <= 2'h0;
    end else if (_T_463) begin
      selArrayWire_1 <= _T_461;
    end
    if (reset) begin
      selArrayWire_0 <= 2'h0;
    end else if (_T_410) begin
      selArrayWire_0 <= _T_408;
    end
    if (reset) begin
      selArrayWire_2 <= 2'h0;
    end else if (_T_516) begin
      selArrayWire_2 <= _T_514;
    end
    if (reset) begin
      selArrayWire_3 <= 2'h0;
    end else if (_T_569) begin
      selArrayWire_3 <= _T_567;
    end
    if (reset) begin
      selArrayWire_4 <= 2'h0;
    end else if (_T_622) begin
      selArrayWire_4 <= _T_620;
    end
    if (reset) begin
      selArrayWire_5 <= 2'h0;
    end else if (_T_675) begin
      selArrayWire_5 <= _T_673;
    end
    if (reset) begin
      selArrayWire_6 <= 2'h0;
    end else if (_T_728) begin
      selArrayWire_6 <= _T_726;
    end
    if (reset) begin
      selArrayWire_7 <= 2'h0;
    end else if (_T_781) begin
      selArrayWire_7 <= _T_779;
    end
    if (reset) begin
      selArrayWire_8 <= 2'h0;
    end else if (_T_834) begin
      selArrayWire_8 <= _T_832;
    end
    if (reset) begin
      selArrayWire_9 <= 2'h0;
    end else if (_T_887) begin
      selArrayWire_9 <= _T_885;
    end
    if (reset) begin
      selArrayWire_10 <= 2'h0;
    end else if (_T_940) begin
      selArrayWire_10 <= _T_938;
    end
    if (reset) begin
      selArrayWire_11 <= 2'h0;
    end else if (_T_993) begin
      selArrayWire_11 <= _T_991;
    end
    if (reset) begin
      selArrayWire_12 <= 2'h0;
    end else if (_T_1046) begin
      selArrayWire_12 <= _T_1044;
    end
    if (reset) begin
      selArrayWire_13 <= 2'h0;
    end else if (_T_1099) begin
      selArrayWire_13 <= _T_1097;
    end
    if (reset) begin
      selArrayWire_14 <= 2'h0;
    end else if (_T_1152) begin
      selArrayWire_14 <= _T_1150;
    end
    if (reset) begin
      selArrayWire_15 <= 2'h0;
    end else if (_T_1205) begin
      selArrayWire_15 <= _T_1203;
    end
    if (reset) begin
      selArrayWire_16 <= 2'h0;
    end else if (_T_1258) begin
      selArrayWire_16 <= _T_1256;
    end
    if (reset) begin
      selArrayWire_17 <= 2'h0;
    end else if (_T_1311) begin
      selArrayWire_17 <= _T_1309;
    end
    if (reset) begin
      selArrayWire_18 <= 2'h0;
    end else if (_T_1364) begin
      selArrayWire_18 <= _T_1362;
    end
    if (reset) begin
      selArrayWire_19 <= 2'h0;
    end else if (_T_1417) begin
      selArrayWire_19 <= _T_1415;
    end
    if (reset) begin
      selArrayWire_20 <= 2'h0;
    end else if (_T_1470) begin
      selArrayWire_20 <= _T_1468;
    end
    if (reset) begin
      selArrayWire_21 <= 2'h0;
    end else if (_T_1523) begin
      selArrayWire_21 <= _T_1521;
    end
    if (reset) begin
      selArrayWire_22 <= 2'h0;
    end else if (_T_1576) begin
      selArrayWire_22 <= _T_1574;
    end
    if (reset) begin
      selArrayWire_23 <= 2'h0;
    end else if (_T_1629) begin
      selArrayWire_23 <= _T_1627;
    end
    if (reset) begin
      selArrayWire_24 <= 2'h0;
    end else if (_T_1682) begin
      selArrayWire_24 <= _T_1680;
    end
    if (reset) begin
      selArrayWire_25 <= 2'h0;
    end else if (_T_1735) begin
      selArrayWire_25 <= _T_1733;
    end
    if (reset) begin
      selArrayWire_26 <= 2'h0;
    end else if (_T_1788) begin
      selArrayWire_26 <= _T_1786;
    end
    if (reset) begin
      selArrayWire_27 <= 2'h0;
    end else if (_T_1841) begin
      selArrayWire_27 <= _T_1839;
    end
    if (reset) begin
      selArrayWire_28 <= 2'h0;
    end else if (_T_1894) begin
      selArrayWire_28 <= _T_1892;
    end
    if (reset) begin
      selArrayWire_29 <= 2'h0;
    end else if (_T_1947) begin
      selArrayWire_29 <= _T_1945;
    end
    if (reset) begin
      selArrayWire_30 <= 2'h0;
    end else if (_T_2000) begin
      selArrayWire_30 <= _T_1998;
    end
    if (reset) begin
      selArrayWire_31 <= 2'h0;
    end else if (_T_2053) begin
      selArrayWire_31 <= _T_2051;
    end
    if (reset) begin
      selArrayWire_32 <= 2'h0;
    end else if (_T_2106) begin
      selArrayWire_32 <= _T_2104;
    end
    if (reset) begin
      selArrayWire_33 <= 2'h0;
    end else if (_T_2159) begin
      selArrayWire_33 <= _T_2157;
    end
    if (reset) begin
      selArrayWire_34 <= 2'h0;
    end else if (_T_2212) begin
      selArrayWire_34 <= _T_2210;
    end
    if (reset) begin
      selArrayWire_35 <= 2'h0;
    end else if (_T_2265) begin
      selArrayWire_35 <= _T_2263;
    end
    if (reset) begin
      selArrayWire_36 <= 2'h0;
    end else if (_T_2318) begin
      selArrayWire_36 <= _T_2316;
    end
    if (reset) begin
      selArrayWire_37 <= 2'h0;
    end else if (_T_2371) begin
      selArrayWire_37 <= _T_2369;
    end
    if (reset) begin
      selArrayWire_38 <= 2'h0;
    end else if (_T_2424) begin
      selArrayWire_38 <= _T_2422;
    end
    if (reset) begin
      selArrayWire_39 <= 2'h0;
    end else if (_T_2477) begin
      selArrayWire_39 <= _T_2475;
    end
    if (reset) begin
      selArrayWire_40 <= 2'h0;
    end else if (_T_2530) begin
      selArrayWire_40 <= _T_2528;
    end
    if (reset) begin
      selArrayWire_41 <= 2'h0;
    end else if (_T_2583) begin
      selArrayWire_41 <= _T_2581;
    end
    if (reset) begin
      selArrayWire_42 <= 2'h0;
    end else if (_T_2636) begin
      selArrayWire_42 <= _T_2634;
    end
    if (reset) begin
      selArrayWire_43 <= 2'h0;
    end else if (_T_2689) begin
      selArrayWire_43 <= _T_2687;
    end
    if (reset) begin
      selArrayWire_44 <= 2'h0;
    end else if (_T_2742) begin
      selArrayWire_44 <= _T_2740;
    end
    if (reset) begin
      selArrayWire_45 <= 2'h0;
    end else if (_T_2795) begin
      selArrayWire_45 <= _T_2793;
    end
    if (reset) begin
      selArrayWire_46 <= 2'h0;
    end else if (_T_2848) begin
      selArrayWire_46 <= _T_2846;
    end
    if (reset) begin
      selArrayWire_47 <= 2'h0;
    end else if (_T_2901) begin
      selArrayWire_47 <= _T_2899;
    end
    if (reset) begin
      selArrayWire_48 <= 2'h0;
    end else if (_T_2954) begin
      selArrayWire_48 <= _T_2952;
    end
    if (reset) begin
      selArrayWire_49 <= 2'h0;
    end else if (_T_3007) begin
      selArrayWire_49 <= _T_3005;
    end
    if (reset) begin
      selArrayWire_50 <= 2'h0;
    end else if (_T_3060) begin
      selArrayWire_50 <= _T_3058;
    end
    if (reset) begin
      selArrayWire_51 <= 2'h0;
    end else if (_T_3113) begin
      selArrayWire_51 <= _T_3111;
    end
    if (reset) begin
      selArrayWire_52 <= 2'h0;
    end else if (_T_3166) begin
      selArrayWire_52 <= _T_3164;
    end
    if (reset) begin
      selArrayWire_53 <= 2'h0;
    end else if (_T_3219) begin
      selArrayWire_53 <= _T_3217;
    end
    if (reset) begin
      selArrayWire_54 <= 2'h0;
    end else if (_T_3272) begin
      selArrayWire_54 <= _T_3270;
    end
    if (reset) begin
      selArrayWire_55 <= 2'h0;
    end else if (_T_3325) begin
      selArrayWire_55 <= _T_3323;
    end
    if (reset) begin
      selArrayWire_56 <= 2'h0;
    end else if (_T_3378) begin
      selArrayWire_56 <= _T_3376;
    end
    if (reset) begin
      selArrayWire_57 <= 2'h0;
    end else if (_T_3431) begin
      selArrayWire_57 <= _T_3429;
    end
    if (reset) begin
      selArrayWire_58 <= 2'h0;
    end else if (_T_3484) begin
      selArrayWire_58 <= _T_3482;
    end
    if (reset) begin
      selArrayWire_59 <= 2'h0;
    end else if (_T_3537) begin
      selArrayWire_59 <= _T_3535;
    end
    if (reset) begin
      selArrayWire_60 <= 2'h0;
    end else if (_T_3590) begin
      selArrayWire_60 <= _T_3588;
    end
    if (reset) begin
      selArrayWire_61 <= 2'h0;
    end else if (_T_3643) begin
      selArrayWire_61 <= _T_3641;
    end
    if (reset) begin
      selArrayWire_62 <= 2'h0;
    end else if (_T_3696) begin
      selArrayWire_62 <= _T_3694;
    end
    if (reset) begin
      selArrayWire_63 <= 2'h0;
    end else if (_T_3749) begin
      selArrayWire_63 <= _T_3747;
    end
  end
endmodule
module clint(
  input         clock,
  input         reset,
  input         io_clintIO_valid,
  output [63:0] io_clintIO_data_read,
  input  [63:0] io_clintIO_data_write,
  input         io_clintIO_wen,
  input  [31:0] io_clintIO_addr,
  output        intrTimeCnt_0,
  input         startTimeCnt_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Reg.scala 27:20]
  wire [63:0] _T_1 = mtime + 64'h1; // @[clint.scala 21:30]
  wire  _T_3 = io_clintIO_valid & io_clintIO_wen; // @[clint.scala 23:70]
  wire  _T_6 = io_clintIO_addr == 32'h2004000; // @[clint.scala 23:105]
  wire  _T_7 = _T_3 & _T_6; // @[clint.scala 23:87]
  reg [63:0] mtimecmp; // @[Reg.scala 27:20]
  wire  _T_13 = 32'h2004000 == io_clintIO_addr; // @[Mux.scala 80:60]
  wire [63:0] _T_14 = _T_13 ? mtimecmp : 64'h0; // @[Mux.scala 80:57]
  wire  _T_15 = 32'h200bff8 == io_clintIO_addr; // @[Mux.scala 80:60]
  wire  _T_17 = mtime >= mtimecmp; // @[clint.scala 37:24]
  wire  _T_18 = _T_17 & startTimeCnt_0; // @[clint.scala 37:36]
  wire  intrTimeCnt = _T_18; // @[clint.scala 36:25 clint.scala 37:15]
  assign io_clintIO_data_read = _T_15 ? mtime : _T_14; // @[clint.scala 27:24]
  assign intrTimeCnt_0 = intrTimeCnt;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mtime <= 64'h0;
    end else if (startTimeCnt_0) begin
      mtime <= _T_1;
    end
    if (reset) begin
      mtimecmp <= 64'h0;
    end else if (_T_7) begin
      mtimecmp <= io_clintIO_data_write;
    end
  end
endmodule
module mem(
  input          clock,
  input          io_memIO_cen,
  input          io_memIO_wen,
  input  [127:0] io_memIO_wdata,
  input  [5:0]   io_memIO_addr,
  input  [127:0] io_memIO_wmask,
  output [127:0] io_memIO_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  cen = ~io_memIO_cen; // @[mem.scala 14:14]
  wire [127:0] bwen = ~io_memIO_wmask; // @[mem.scala 15:15]
  wire  wen = ~io_memIO_wen; // @[mem.scala 16:14]
  wire [127:0] _T_2 = io_memIO_wdata & bwen; // @[mem.scala 25:47]
  reg [127:0] ramWire_0; // @[Reg.scala 15:16]
  wire [127:0] _T_3 = ramWire_0 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_4 = _T_2 | _T_3; // @[mem.scala 25:55]
  wire  _T_5 = cen & wen; // @[mem.scala 25:91]
  wire  _T_6 = io_memIO_addr == 6'h0; // @[mem.scala 25:115]
  wire  _T_7 = _T_5 & _T_6; // @[mem.scala 25:98]
  reg [127:0] ramWire_1; // @[Reg.scala 15:16]
  wire [127:0] _T_10 = ramWire_1 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_11 = _T_2 | _T_10; // @[mem.scala 25:55]
  wire  _T_13 = io_memIO_addr == 6'h1; // @[mem.scala 25:115]
  wire  _T_14 = _T_5 & _T_13; // @[mem.scala 25:98]
  reg [127:0] ramWire_2; // @[Reg.scala 15:16]
  wire [127:0] _T_17 = ramWire_2 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_18 = _T_2 | _T_17; // @[mem.scala 25:55]
  wire  _T_20 = io_memIO_addr == 6'h2; // @[mem.scala 25:115]
  wire  _T_21 = _T_5 & _T_20; // @[mem.scala 25:98]
  reg [127:0] ramWire_3; // @[Reg.scala 15:16]
  wire [127:0] _T_24 = ramWire_3 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_25 = _T_2 | _T_24; // @[mem.scala 25:55]
  wire  _T_27 = io_memIO_addr == 6'h3; // @[mem.scala 25:115]
  wire  _T_28 = _T_5 & _T_27; // @[mem.scala 25:98]
  reg [127:0] ramWire_4; // @[Reg.scala 15:16]
  wire [127:0] _T_31 = ramWire_4 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_32 = _T_2 | _T_31; // @[mem.scala 25:55]
  wire  _T_34 = io_memIO_addr == 6'h4; // @[mem.scala 25:115]
  wire  _T_35 = _T_5 & _T_34; // @[mem.scala 25:98]
  reg [127:0] ramWire_5; // @[Reg.scala 15:16]
  wire [127:0] _T_38 = ramWire_5 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_39 = _T_2 | _T_38; // @[mem.scala 25:55]
  wire  _T_41 = io_memIO_addr == 6'h5; // @[mem.scala 25:115]
  wire  _T_42 = _T_5 & _T_41; // @[mem.scala 25:98]
  reg [127:0] ramWire_6; // @[Reg.scala 15:16]
  wire [127:0] _T_45 = ramWire_6 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_46 = _T_2 | _T_45; // @[mem.scala 25:55]
  wire  _T_48 = io_memIO_addr == 6'h6; // @[mem.scala 25:115]
  wire  _T_49 = _T_5 & _T_48; // @[mem.scala 25:98]
  reg [127:0] ramWire_7; // @[Reg.scala 15:16]
  wire [127:0] _T_52 = ramWire_7 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_53 = _T_2 | _T_52; // @[mem.scala 25:55]
  wire  _T_55 = io_memIO_addr == 6'h7; // @[mem.scala 25:115]
  wire  _T_56 = _T_5 & _T_55; // @[mem.scala 25:98]
  reg [127:0] ramWire_8; // @[Reg.scala 15:16]
  wire [127:0] _T_59 = ramWire_8 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_60 = _T_2 | _T_59; // @[mem.scala 25:55]
  wire  _T_62 = io_memIO_addr == 6'h8; // @[mem.scala 25:115]
  wire  _T_63 = _T_5 & _T_62; // @[mem.scala 25:98]
  reg [127:0] ramWire_9; // @[Reg.scala 15:16]
  wire [127:0] _T_66 = ramWire_9 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_67 = _T_2 | _T_66; // @[mem.scala 25:55]
  wire  _T_69 = io_memIO_addr == 6'h9; // @[mem.scala 25:115]
  wire  _T_70 = _T_5 & _T_69; // @[mem.scala 25:98]
  reg [127:0] ramWire_10; // @[Reg.scala 15:16]
  wire [127:0] _T_73 = ramWire_10 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_74 = _T_2 | _T_73; // @[mem.scala 25:55]
  wire  _T_76 = io_memIO_addr == 6'ha; // @[mem.scala 25:115]
  wire  _T_77 = _T_5 & _T_76; // @[mem.scala 25:98]
  reg [127:0] ramWire_11; // @[Reg.scala 15:16]
  wire [127:0] _T_80 = ramWire_11 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_81 = _T_2 | _T_80; // @[mem.scala 25:55]
  wire  _T_83 = io_memIO_addr == 6'hb; // @[mem.scala 25:115]
  wire  _T_84 = _T_5 & _T_83; // @[mem.scala 25:98]
  reg [127:0] ramWire_12; // @[Reg.scala 15:16]
  wire [127:0] _T_87 = ramWire_12 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_88 = _T_2 | _T_87; // @[mem.scala 25:55]
  wire  _T_90 = io_memIO_addr == 6'hc; // @[mem.scala 25:115]
  wire  _T_91 = _T_5 & _T_90; // @[mem.scala 25:98]
  reg [127:0] ramWire_13; // @[Reg.scala 15:16]
  wire [127:0] _T_94 = ramWire_13 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_95 = _T_2 | _T_94; // @[mem.scala 25:55]
  wire  _T_97 = io_memIO_addr == 6'hd; // @[mem.scala 25:115]
  wire  _T_98 = _T_5 & _T_97; // @[mem.scala 25:98]
  reg [127:0] ramWire_14; // @[Reg.scala 15:16]
  wire [127:0] _T_101 = ramWire_14 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_102 = _T_2 | _T_101; // @[mem.scala 25:55]
  wire  _T_104 = io_memIO_addr == 6'he; // @[mem.scala 25:115]
  wire  _T_105 = _T_5 & _T_104; // @[mem.scala 25:98]
  reg [127:0] ramWire_15; // @[Reg.scala 15:16]
  wire [127:0] _T_108 = ramWire_15 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_109 = _T_2 | _T_108; // @[mem.scala 25:55]
  wire  _T_111 = io_memIO_addr == 6'hf; // @[mem.scala 25:115]
  wire  _T_112 = _T_5 & _T_111; // @[mem.scala 25:98]
  reg [127:0] ramWire_16; // @[Reg.scala 15:16]
  wire [127:0] _T_115 = ramWire_16 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_116 = _T_2 | _T_115; // @[mem.scala 25:55]
  wire  _T_118 = io_memIO_addr == 6'h10; // @[mem.scala 25:115]
  wire  _T_119 = _T_5 & _T_118; // @[mem.scala 25:98]
  reg [127:0] ramWire_17; // @[Reg.scala 15:16]
  wire [127:0] _T_122 = ramWire_17 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_123 = _T_2 | _T_122; // @[mem.scala 25:55]
  wire  _T_125 = io_memIO_addr == 6'h11; // @[mem.scala 25:115]
  wire  _T_126 = _T_5 & _T_125; // @[mem.scala 25:98]
  reg [127:0] ramWire_18; // @[Reg.scala 15:16]
  wire [127:0] _T_129 = ramWire_18 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_130 = _T_2 | _T_129; // @[mem.scala 25:55]
  wire  _T_132 = io_memIO_addr == 6'h12; // @[mem.scala 25:115]
  wire  _T_133 = _T_5 & _T_132; // @[mem.scala 25:98]
  reg [127:0] ramWire_19; // @[Reg.scala 15:16]
  wire [127:0] _T_136 = ramWire_19 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_137 = _T_2 | _T_136; // @[mem.scala 25:55]
  wire  _T_139 = io_memIO_addr == 6'h13; // @[mem.scala 25:115]
  wire  _T_140 = _T_5 & _T_139; // @[mem.scala 25:98]
  reg [127:0] ramWire_20; // @[Reg.scala 15:16]
  wire [127:0] _T_143 = ramWire_20 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_144 = _T_2 | _T_143; // @[mem.scala 25:55]
  wire  _T_146 = io_memIO_addr == 6'h14; // @[mem.scala 25:115]
  wire  _T_147 = _T_5 & _T_146; // @[mem.scala 25:98]
  reg [127:0] ramWire_21; // @[Reg.scala 15:16]
  wire [127:0] _T_150 = ramWire_21 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_151 = _T_2 | _T_150; // @[mem.scala 25:55]
  wire  _T_153 = io_memIO_addr == 6'h15; // @[mem.scala 25:115]
  wire  _T_154 = _T_5 & _T_153; // @[mem.scala 25:98]
  reg [127:0] ramWire_22; // @[Reg.scala 15:16]
  wire [127:0] _T_157 = ramWire_22 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_158 = _T_2 | _T_157; // @[mem.scala 25:55]
  wire  _T_160 = io_memIO_addr == 6'h16; // @[mem.scala 25:115]
  wire  _T_161 = _T_5 & _T_160; // @[mem.scala 25:98]
  reg [127:0] ramWire_23; // @[Reg.scala 15:16]
  wire [127:0] _T_164 = ramWire_23 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_165 = _T_2 | _T_164; // @[mem.scala 25:55]
  wire  _T_167 = io_memIO_addr == 6'h17; // @[mem.scala 25:115]
  wire  _T_168 = _T_5 & _T_167; // @[mem.scala 25:98]
  reg [127:0] ramWire_24; // @[Reg.scala 15:16]
  wire [127:0] _T_171 = ramWire_24 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_172 = _T_2 | _T_171; // @[mem.scala 25:55]
  wire  _T_174 = io_memIO_addr == 6'h18; // @[mem.scala 25:115]
  wire  _T_175 = _T_5 & _T_174; // @[mem.scala 25:98]
  reg [127:0] ramWire_25; // @[Reg.scala 15:16]
  wire [127:0] _T_178 = ramWire_25 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_179 = _T_2 | _T_178; // @[mem.scala 25:55]
  wire  _T_181 = io_memIO_addr == 6'h19; // @[mem.scala 25:115]
  wire  _T_182 = _T_5 & _T_181; // @[mem.scala 25:98]
  reg [127:0] ramWire_26; // @[Reg.scala 15:16]
  wire [127:0] _T_185 = ramWire_26 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_186 = _T_2 | _T_185; // @[mem.scala 25:55]
  wire  _T_188 = io_memIO_addr == 6'h1a; // @[mem.scala 25:115]
  wire  _T_189 = _T_5 & _T_188; // @[mem.scala 25:98]
  reg [127:0] ramWire_27; // @[Reg.scala 15:16]
  wire [127:0] _T_192 = ramWire_27 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_193 = _T_2 | _T_192; // @[mem.scala 25:55]
  wire  _T_195 = io_memIO_addr == 6'h1b; // @[mem.scala 25:115]
  wire  _T_196 = _T_5 & _T_195; // @[mem.scala 25:98]
  reg [127:0] ramWire_28; // @[Reg.scala 15:16]
  wire [127:0] _T_199 = ramWire_28 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_200 = _T_2 | _T_199; // @[mem.scala 25:55]
  wire  _T_202 = io_memIO_addr == 6'h1c; // @[mem.scala 25:115]
  wire  _T_203 = _T_5 & _T_202; // @[mem.scala 25:98]
  reg [127:0] ramWire_29; // @[Reg.scala 15:16]
  wire [127:0] _T_206 = ramWire_29 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_207 = _T_2 | _T_206; // @[mem.scala 25:55]
  wire  _T_209 = io_memIO_addr == 6'h1d; // @[mem.scala 25:115]
  wire  _T_210 = _T_5 & _T_209; // @[mem.scala 25:98]
  reg [127:0] ramWire_30; // @[Reg.scala 15:16]
  wire [127:0] _T_213 = ramWire_30 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_214 = _T_2 | _T_213; // @[mem.scala 25:55]
  wire  _T_216 = io_memIO_addr == 6'h1e; // @[mem.scala 25:115]
  wire  _T_217 = _T_5 & _T_216; // @[mem.scala 25:98]
  reg [127:0] ramWire_31; // @[Reg.scala 15:16]
  wire [127:0] _T_220 = ramWire_31 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_221 = _T_2 | _T_220; // @[mem.scala 25:55]
  wire  _T_223 = io_memIO_addr == 6'h1f; // @[mem.scala 25:115]
  wire  _T_224 = _T_5 & _T_223; // @[mem.scala 25:98]
  reg [127:0] ramWire_32; // @[Reg.scala 15:16]
  wire [127:0] _T_227 = ramWire_32 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_228 = _T_2 | _T_227; // @[mem.scala 25:55]
  wire  _T_230 = io_memIO_addr == 6'h20; // @[mem.scala 25:115]
  wire  _T_231 = _T_5 & _T_230; // @[mem.scala 25:98]
  reg [127:0] ramWire_33; // @[Reg.scala 15:16]
  wire [127:0] _T_234 = ramWire_33 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_235 = _T_2 | _T_234; // @[mem.scala 25:55]
  wire  _T_237 = io_memIO_addr == 6'h21; // @[mem.scala 25:115]
  wire  _T_238 = _T_5 & _T_237; // @[mem.scala 25:98]
  reg [127:0] ramWire_34; // @[Reg.scala 15:16]
  wire [127:0] _T_241 = ramWire_34 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_242 = _T_2 | _T_241; // @[mem.scala 25:55]
  wire  _T_244 = io_memIO_addr == 6'h22; // @[mem.scala 25:115]
  wire  _T_245 = _T_5 & _T_244; // @[mem.scala 25:98]
  reg [127:0] ramWire_35; // @[Reg.scala 15:16]
  wire [127:0] _T_248 = ramWire_35 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_249 = _T_2 | _T_248; // @[mem.scala 25:55]
  wire  _T_251 = io_memIO_addr == 6'h23; // @[mem.scala 25:115]
  wire  _T_252 = _T_5 & _T_251; // @[mem.scala 25:98]
  reg [127:0] ramWire_36; // @[Reg.scala 15:16]
  wire [127:0] _T_255 = ramWire_36 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_256 = _T_2 | _T_255; // @[mem.scala 25:55]
  wire  _T_258 = io_memIO_addr == 6'h24; // @[mem.scala 25:115]
  wire  _T_259 = _T_5 & _T_258; // @[mem.scala 25:98]
  reg [127:0] ramWire_37; // @[Reg.scala 15:16]
  wire [127:0] _T_262 = ramWire_37 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_263 = _T_2 | _T_262; // @[mem.scala 25:55]
  wire  _T_265 = io_memIO_addr == 6'h25; // @[mem.scala 25:115]
  wire  _T_266 = _T_5 & _T_265; // @[mem.scala 25:98]
  reg [127:0] ramWire_38; // @[Reg.scala 15:16]
  wire [127:0] _T_269 = ramWire_38 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_270 = _T_2 | _T_269; // @[mem.scala 25:55]
  wire  _T_272 = io_memIO_addr == 6'h26; // @[mem.scala 25:115]
  wire  _T_273 = _T_5 & _T_272; // @[mem.scala 25:98]
  reg [127:0] ramWire_39; // @[Reg.scala 15:16]
  wire [127:0] _T_276 = ramWire_39 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_277 = _T_2 | _T_276; // @[mem.scala 25:55]
  wire  _T_279 = io_memIO_addr == 6'h27; // @[mem.scala 25:115]
  wire  _T_280 = _T_5 & _T_279; // @[mem.scala 25:98]
  reg [127:0] ramWire_40; // @[Reg.scala 15:16]
  wire [127:0] _T_283 = ramWire_40 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_284 = _T_2 | _T_283; // @[mem.scala 25:55]
  wire  _T_286 = io_memIO_addr == 6'h28; // @[mem.scala 25:115]
  wire  _T_287 = _T_5 & _T_286; // @[mem.scala 25:98]
  reg [127:0] ramWire_41; // @[Reg.scala 15:16]
  wire [127:0] _T_290 = ramWire_41 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_291 = _T_2 | _T_290; // @[mem.scala 25:55]
  wire  _T_293 = io_memIO_addr == 6'h29; // @[mem.scala 25:115]
  wire  _T_294 = _T_5 & _T_293; // @[mem.scala 25:98]
  reg [127:0] ramWire_42; // @[Reg.scala 15:16]
  wire [127:0] _T_297 = ramWire_42 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_298 = _T_2 | _T_297; // @[mem.scala 25:55]
  wire  _T_300 = io_memIO_addr == 6'h2a; // @[mem.scala 25:115]
  wire  _T_301 = _T_5 & _T_300; // @[mem.scala 25:98]
  reg [127:0] ramWire_43; // @[Reg.scala 15:16]
  wire [127:0] _T_304 = ramWire_43 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_305 = _T_2 | _T_304; // @[mem.scala 25:55]
  wire  _T_307 = io_memIO_addr == 6'h2b; // @[mem.scala 25:115]
  wire  _T_308 = _T_5 & _T_307; // @[mem.scala 25:98]
  reg [127:0] ramWire_44; // @[Reg.scala 15:16]
  wire [127:0] _T_311 = ramWire_44 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_312 = _T_2 | _T_311; // @[mem.scala 25:55]
  wire  _T_314 = io_memIO_addr == 6'h2c; // @[mem.scala 25:115]
  wire  _T_315 = _T_5 & _T_314; // @[mem.scala 25:98]
  reg [127:0] ramWire_45; // @[Reg.scala 15:16]
  wire [127:0] _T_318 = ramWire_45 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_319 = _T_2 | _T_318; // @[mem.scala 25:55]
  wire  _T_321 = io_memIO_addr == 6'h2d; // @[mem.scala 25:115]
  wire  _T_322 = _T_5 & _T_321; // @[mem.scala 25:98]
  reg [127:0] ramWire_46; // @[Reg.scala 15:16]
  wire [127:0] _T_325 = ramWire_46 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_326 = _T_2 | _T_325; // @[mem.scala 25:55]
  wire  _T_328 = io_memIO_addr == 6'h2e; // @[mem.scala 25:115]
  wire  _T_329 = _T_5 & _T_328; // @[mem.scala 25:98]
  reg [127:0] ramWire_47; // @[Reg.scala 15:16]
  wire [127:0] _T_332 = ramWire_47 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_333 = _T_2 | _T_332; // @[mem.scala 25:55]
  wire  _T_335 = io_memIO_addr == 6'h2f; // @[mem.scala 25:115]
  wire  _T_336 = _T_5 & _T_335; // @[mem.scala 25:98]
  reg [127:0] ramWire_48; // @[Reg.scala 15:16]
  wire [127:0] _T_339 = ramWire_48 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_340 = _T_2 | _T_339; // @[mem.scala 25:55]
  wire  _T_342 = io_memIO_addr == 6'h30; // @[mem.scala 25:115]
  wire  _T_343 = _T_5 & _T_342; // @[mem.scala 25:98]
  reg [127:0] ramWire_49; // @[Reg.scala 15:16]
  wire [127:0] _T_346 = ramWire_49 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_347 = _T_2 | _T_346; // @[mem.scala 25:55]
  wire  _T_349 = io_memIO_addr == 6'h31; // @[mem.scala 25:115]
  wire  _T_350 = _T_5 & _T_349; // @[mem.scala 25:98]
  reg [127:0] ramWire_50; // @[Reg.scala 15:16]
  wire [127:0] _T_353 = ramWire_50 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_354 = _T_2 | _T_353; // @[mem.scala 25:55]
  wire  _T_356 = io_memIO_addr == 6'h32; // @[mem.scala 25:115]
  wire  _T_357 = _T_5 & _T_356; // @[mem.scala 25:98]
  reg [127:0] ramWire_51; // @[Reg.scala 15:16]
  wire [127:0] _T_360 = ramWire_51 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_361 = _T_2 | _T_360; // @[mem.scala 25:55]
  wire  _T_363 = io_memIO_addr == 6'h33; // @[mem.scala 25:115]
  wire  _T_364 = _T_5 & _T_363; // @[mem.scala 25:98]
  reg [127:0] ramWire_52; // @[Reg.scala 15:16]
  wire [127:0] _T_367 = ramWire_52 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_368 = _T_2 | _T_367; // @[mem.scala 25:55]
  wire  _T_370 = io_memIO_addr == 6'h34; // @[mem.scala 25:115]
  wire  _T_371 = _T_5 & _T_370; // @[mem.scala 25:98]
  reg [127:0] ramWire_53; // @[Reg.scala 15:16]
  wire [127:0] _T_374 = ramWire_53 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_375 = _T_2 | _T_374; // @[mem.scala 25:55]
  wire  _T_377 = io_memIO_addr == 6'h35; // @[mem.scala 25:115]
  wire  _T_378 = _T_5 & _T_377; // @[mem.scala 25:98]
  reg [127:0] ramWire_54; // @[Reg.scala 15:16]
  wire [127:0] _T_381 = ramWire_54 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_382 = _T_2 | _T_381; // @[mem.scala 25:55]
  wire  _T_384 = io_memIO_addr == 6'h36; // @[mem.scala 25:115]
  wire  _T_385 = _T_5 & _T_384; // @[mem.scala 25:98]
  reg [127:0] ramWire_55; // @[Reg.scala 15:16]
  wire [127:0] _T_388 = ramWire_55 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_389 = _T_2 | _T_388; // @[mem.scala 25:55]
  wire  _T_391 = io_memIO_addr == 6'h37; // @[mem.scala 25:115]
  wire  _T_392 = _T_5 & _T_391; // @[mem.scala 25:98]
  reg [127:0] ramWire_56; // @[Reg.scala 15:16]
  wire [127:0] _T_395 = ramWire_56 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_396 = _T_2 | _T_395; // @[mem.scala 25:55]
  wire  _T_398 = io_memIO_addr == 6'h38; // @[mem.scala 25:115]
  wire  _T_399 = _T_5 & _T_398; // @[mem.scala 25:98]
  reg [127:0] ramWire_57; // @[Reg.scala 15:16]
  wire [127:0] _T_402 = ramWire_57 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_403 = _T_2 | _T_402; // @[mem.scala 25:55]
  wire  _T_405 = io_memIO_addr == 6'h39; // @[mem.scala 25:115]
  wire  _T_406 = _T_5 & _T_405; // @[mem.scala 25:98]
  reg [127:0] ramWire_58; // @[Reg.scala 15:16]
  wire [127:0] _T_409 = ramWire_58 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_410 = _T_2 | _T_409; // @[mem.scala 25:55]
  wire  _T_412 = io_memIO_addr == 6'h3a; // @[mem.scala 25:115]
  wire  _T_413 = _T_5 & _T_412; // @[mem.scala 25:98]
  reg [127:0] ramWire_59; // @[Reg.scala 15:16]
  wire [127:0] _T_416 = ramWire_59 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_417 = _T_2 | _T_416; // @[mem.scala 25:55]
  wire  _T_419 = io_memIO_addr == 6'h3b; // @[mem.scala 25:115]
  wire  _T_420 = _T_5 & _T_419; // @[mem.scala 25:98]
  reg [127:0] ramWire_60; // @[Reg.scala 15:16]
  wire [127:0] _T_423 = ramWire_60 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_424 = _T_2 | _T_423; // @[mem.scala 25:55]
  wire  _T_426 = io_memIO_addr == 6'h3c; // @[mem.scala 25:115]
  wire  _T_427 = _T_5 & _T_426; // @[mem.scala 25:98]
  reg [127:0] ramWire_61; // @[Reg.scala 15:16]
  wire [127:0] _T_430 = ramWire_61 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_431 = _T_2 | _T_430; // @[mem.scala 25:55]
  wire  _T_433 = io_memIO_addr == 6'h3d; // @[mem.scala 25:115]
  wire  _T_434 = _T_5 & _T_433; // @[mem.scala 25:98]
  reg [127:0] ramWire_62; // @[Reg.scala 15:16]
  wire [127:0] _T_437 = ramWire_62 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_438 = _T_2 | _T_437; // @[mem.scala 25:55]
  wire  _T_440 = io_memIO_addr == 6'h3e; // @[mem.scala 25:115]
  wire  _T_441 = _T_5 & _T_440; // @[mem.scala 25:98]
  reg [127:0] ramWire_63; // @[Reg.scala 15:16]
  wire [127:0] _T_444 = ramWire_63 & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _T_445 = _T_2 | _T_444; // @[mem.scala 25:55]
  wire  _T_447 = io_memIO_addr == 6'h3f; // @[mem.scala 25:115]
  wire  _T_448 = _T_5 & _T_447; // @[mem.scala 25:98]
  wire  _T_450 = 6'h1 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_451 = _T_450 ? ramWire_1 : ramWire_0; // @[Mux.scala 80:57]
  wire  _T_452 = 6'h2 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_453 = _T_452 ? ramWire_2 : _T_451; // @[Mux.scala 80:57]
  wire  _T_454 = 6'h3 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_455 = _T_454 ? ramWire_3 : _T_453; // @[Mux.scala 80:57]
  wire  _T_456 = 6'h4 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_457 = _T_456 ? ramWire_4 : _T_455; // @[Mux.scala 80:57]
  wire  _T_458 = 6'h5 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_459 = _T_458 ? ramWire_5 : _T_457; // @[Mux.scala 80:57]
  wire  _T_460 = 6'h6 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_461 = _T_460 ? ramWire_6 : _T_459; // @[Mux.scala 80:57]
  wire  _T_462 = 6'h7 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_463 = _T_462 ? ramWire_7 : _T_461; // @[Mux.scala 80:57]
  wire  _T_464 = 6'h8 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_465 = _T_464 ? ramWire_8 : _T_463; // @[Mux.scala 80:57]
  wire  _T_466 = 6'h9 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_467 = _T_466 ? ramWire_9 : _T_465; // @[Mux.scala 80:57]
  wire  _T_468 = 6'ha == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_469 = _T_468 ? ramWire_10 : _T_467; // @[Mux.scala 80:57]
  wire  _T_470 = 6'hb == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_471 = _T_470 ? ramWire_11 : _T_469; // @[Mux.scala 80:57]
  wire  _T_472 = 6'hc == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_473 = _T_472 ? ramWire_12 : _T_471; // @[Mux.scala 80:57]
  wire  _T_474 = 6'hd == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_475 = _T_474 ? ramWire_13 : _T_473; // @[Mux.scala 80:57]
  wire  _T_476 = 6'he == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_477 = _T_476 ? ramWire_14 : _T_475; // @[Mux.scala 80:57]
  wire  _T_478 = 6'hf == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_479 = _T_478 ? ramWire_15 : _T_477; // @[Mux.scala 80:57]
  wire  _T_480 = 6'h10 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_481 = _T_480 ? ramWire_16 : _T_479; // @[Mux.scala 80:57]
  wire  _T_482 = 6'h11 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_483 = _T_482 ? ramWire_17 : _T_481; // @[Mux.scala 80:57]
  wire  _T_484 = 6'h12 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_485 = _T_484 ? ramWire_18 : _T_483; // @[Mux.scala 80:57]
  wire  _T_486 = 6'h13 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_487 = _T_486 ? ramWire_19 : _T_485; // @[Mux.scala 80:57]
  wire  _T_488 = 6'h14 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_489 = _T_488 ? ramWire_20 : _T_487; // @[Mux.scala 80:57]
  wire  _T_490 = 6'h15 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_491 = _T_490 ? ramWire_21 : _T_489; // @[Mux.scala 80:57]
  wire  _T_492 = 6'h16 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_493 = _T_492 ? ramWire_22 : _T_491; // @[Mux.scala 80:57]
  wire  _T_494 = 6'h17 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_495 = _T_494 ? ramWire_23 : _T_493; // @[Mux.scala 80:57]
  wire  _T_496 = 6'h18 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_497 = _T_496 ? ramWire_24 : _T_495; // @[Mux.scala 80:57]
  wire  _T_498 = 6'h19 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_499 = _T_498 ? ramWire_25 : _T_497; // @[Mux.scala 80:57]
  wire  _T_500 = 6'h1a == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_501 = _T_500 ? ramWire_26 : _T_499; // @[Mux.scala 80:57]
  wire  _T_502 = 6'h1b == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_503 = _T_502 ? ramWire_27 : _T_501; // @[Mux.scala 80:57]
  wire  _T_504 = 6'h1c == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_505 = _T_504 ? ramWire_28 : _T_503; // @[Mux.scala 80:57]
  wire  _T_506 = 6'h1d == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_507 = _T_506 ? ramWire_29 : _T_505; // @[Mux.scala 80:57]
  wire  _T_508 = 6'h1e == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_509 = _T_508 ? ramWire_30 : _T_507; // @[Mux.scala 80:57]
  wire  _T_510 = 6'h1f == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_511 = _T_510 ? ramWire_31 : _T_509; // @[Mux.scala 80:57]
  wire  _T_512 = 6'h20 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_513 = _T_512 ? ramWire_32 : _T_511; // @[Mux.scala 80:57]
  wire  _T_514 = 6'h21 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_515 = _T_514 ? ramWire_33 : _T_513; // @[Mux.scala 80:57]
  wire  _T_516 = 6'h22 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_517 = _T_516 ? ramWire_34 : _T_515; // @[Mux.scala 80:57]
  wire  _T_518 = 6'h23 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_519 = _T_518 ? ramWire_35 : _T_517; // @[Mux.scala 80:57]
  wire  _T_520 = 6'h24 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_521 = _T_520 ? ramWire_36 : _T_519; // @[Mux.scala 80:57]
  wire  _T_522 = 6'h25 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_523 = _T_522 ? ramWire_37 : _T_521; // @[Mux.scala 80:57]
  wire  _T_524 = 6'h26 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_525 = _T_524 ? ramWire_38 : _T_523; // @[Mux.scala 80:57]
  wire  _T_526 = 6'h27 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_527 = _T_526 ? ramWire_39 : _T_525; // @[Mux.scala 80:57]
  wire  _T_528 = 6'h28 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_529 = _T_528 ? ramWire_40 : _T_527; // @[Mux.scala 80:57]
  wire  _T_530 = 6'h29 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_531 = _T_530 ? ramWire_41 : _T_529; // @[Mux.scala 80:57]
  wire  _T_532 = 6'h2a == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_533 = _T_532 ? ramWire_42 : _T_531; // @[Mux.scala 80:57]
  wire  _T_534 = 6'h2b == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_535 = _T_534 ? ramWire_43 : _T_533; // @[Mux.scala 80:57]
  wire  _T_536 = 6'h2c == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_537 = _T_536 ? ramWire_44 : _T_535; // @[Mux.scala 80:57]
  wire  _T_538 = 6'h2d == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_539 = _T_538 ? ramWire_45 : _T_537; // @[Mux.scala 80:57]
  wire  _T_540 = 6'h2e == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_541 = _T_540 ? ramWire_46 : _T_539; // @[Mux.scala 80:57]
  wire  _T_542 = 6'h2f == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_543 = _T_542 ? ramWire_47 : _T_541; // @[Mux.scala 80:57]
  wire  _T_544 = 6'h30 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_545 = _T_544 ? ramWire_48 : _T_543; // @[Mux.scala 80:57]
  wire  _T_546 = 6'h31 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_547 = _T_546 ? ramWire_49 : _T_545; // @[Mux.scala 80:57]
  wire  _T_548 = 6'h32 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_549 = _T_548 ? ramWire_50 : _T_547; // @[Mux.scala 80:57]
  wire  _T_550 = 6'h33 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_551 = _T_550 ? ramWire_51 : _T_549; // @[Mux.scala 80:57]
  wire  _T_552 = 6'h34 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_553 = _T_552 ? ramWire_52 : _T_551; // @[Mux.scala 80:57]
  wire  _T_554 = 6'h35 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_555 = _T_554 ? ramWire_53 : _T_553; // @[Mux.scala 80:57]
  wire  _T_556 = 6'h36 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_557 = _T_556 ? ramWire_54 : _T_555; // @[Mux.scala 80:57]
  wire  _T_558 = 6'h37 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_559 = _T_558 ? ramWire_55 : _T_557; // @[Mux.scala 80:57]
  wire  _T_560 = 6'h38 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_561 = _T_560 ? ramWire_56 : _T_559; // @[Mux.scala 80:57]
  wire  _T_562 = 6'h39 == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_563 = _T_562 ? ramWire_57 : _T_561; // @[Mux.scala 80:57]
  wire  _T_564 = 6'h3a == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_565 = _T_564 ? ramWire_58 : _T_563; // @[Mux.scala 80:57]
  wire  _T_566 = 6'h3b == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_567 = _T_566 ? ramWire_59 : _T_565; // @[Mux.scala 80:57]
  wire  _T_568 = 6'h3c == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_569 = _T_568 ? ramWire_60 : _T_567; // @[Mux.scala 80:57]
  wire  _T_570 = 6'h3d == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_571 = _T_570 ? ramWire_61 : _T_569; // @[Mux.scala 80:57]
  wire  _T_572 = 6'h3e == io_memIO_addr; // @[Mux.scala 80:60]
  wire [127:0] _T_573 = _T_572 ? ramWire_62 : _T_571; // @[Mux.scala 80:57]
  wire  _T_574 = 6'h3f == io_memIO_addr; // @[Mux.scala 80:60]
  assign io_memIO_rdata = _T_574 ? ramWire_63 : _T_573; // @[mem.scala 30:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  ramWire_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  ramWire_1 = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  ramWire_2 = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  ramWire_3 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  ramWire_4 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  ramWire_5 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  ramWire_6 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  ramWire_7 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  ramWire_8 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  ramWire_9 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  ramWire_10 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  ramWire_11 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  ramWire_12 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  ramWire_13 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  ramWire_14 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  ramWire_15 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  ramWire_16 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  ramWire_17 = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  ramWire_18 = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  ramWire_19 = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  ramWire_20 = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  ramWire_21 = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  ramWire_22 = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  ramWire_23 = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  ramWire_24 = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  ramWire_25 = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  ramWire_26 = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  ramWire_27 = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  ramWire_28 = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  ramWire_29 = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  ramWire_30 = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  ramWire_31 = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  ramWire_32 = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  ramWire_33 = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  ramWire_34 = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  ramWire_35 = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  ramWire_36 = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  ramWire_37 = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  ramWire_38 = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  ramWire_39 = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  ramWire_40 = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  ramWire_41 = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  ramWire_42 = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  ramWire_43 = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  ramWire_44 = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  ramWire_45 = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  ramWire_46 = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  ramWire_47 = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  ramWire_48 = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  ramWire_49 = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  ramWire_50 = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  ramWire_51 = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  ramWire_52 = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  ramWire_53 = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  ramWire_54 = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  ramWire_55 = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  ramWire_56 = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  ramWire_57 = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  ramWire_58 = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  ramWire_59 = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  ramWire_60 = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  ramWire_61 = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  ramWire_62 = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  ramWire_63 = _RAND_63[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_7) begin
      ramWire_0 <= _T_4;
    end
    if (_T_14) begin
      ramWire_1 <= _T_11;
    end
    if (_T_21) begin
      ramWire_2 <= _T_18;
    end
    if (_T_28) begin
      ramWire_3 <= _T_25;
    end
    if (_T_35) begin
      ramWire_4 <= _T_32;
    end
    if (_T_42) begin
      ramWire_5 <= _T_39;
    end
    if (_T_49) begin
      ramWire_6 <= _T_46;
    end
    if (_T_56) begin
      ramWire_7 <= _T_53;
    end
    if (_T_63) begin
      ramWire_8 <= _T_60;
    end
    if (_T_70) begin
      ramWire_9 <= _T_67;
    end
    if (_T_77) begin
      ramWire_10 <= _T_74;
    end
    if (_T_84) begin
      ramWire_11 <= _T_81;
    end
    if (_T_91) begin
      ramWire_12 <= _T_88;
    end
    if (_T_98) begin
      ramWire_13 <= _T_95;
    end
    if (_T_105) begin
      ramWire_14 <= _T_102;
    end
    if (_T_112) begin
      ramWire_15 <= _T_109;
    end
    if (_T_119) begin
      ramWire_16 <= _T_116;
    end
    if (_T_126) begin
      ramWire_17 <= _T_123;
    end
    if (_T_133) begin
      ramWire_18 <= _T_130;
    end
    if (_T_140) begin
      ramWire_19 <= _T_137;
    end
    if (_T_147) begin
      ramWire_20 <= _T_144;
    end
    if (_T_154) begin
      ramWire_21 <= _T_151;
    end
    if (_T_161) begin
      ramWire_22 <= _T_158;
    end
    if (_T_168) begin
      ramWire_23 <= _T_165;
    end
    if (_T_175) begin
      ramWire_24 <= _T_172;
    end
    if (_T_182) begin
      ramWire_25 <= _T_179;
    end
    if (_T_189) begin
      ramWire_26 <= _T_186;
    end
    if (_T_196) begin
      ramWire_27 <= _T_193;
    end
    if (_T_203) begin
      ramWire_28 <= _T_200;
    end
    if (_T_210) begin
      ramWire_29 <= _T_207;
    end
    if (_T_217) begin
      ramWire_30 <= _T_214;
    end
    if (_T_224) begin
      ramWire_31 <= _T_221;
    end
    if (_T_231) begin
      ramWire_32 <= _T_228;
    end
    if (_T_238) begin
      ramWire_33 <= _T_235;
    end
    if (_T_245) begin
      ramWire_34 <= _T_242;
    end
    if (_T_252) begin
      ramWire_35 <= _T_249;
    end
    if (_T_259) begin
      ramWire_36 <= _T_256;
    end
    if (_T_266) begin
      ramWire_37 <= _T_263;
    end
    if (_T_273) begin
      ramWire_38 <= _T_270;
    end
    if (_T_280) begin
      ramWire_39 <= _T_277;
    end
    if (_T_287) begin
      ramWire_40 <= _T_284;
    end
    if (_T_294) begin
      ramWire_41 <= _T_291;
    end
    if (_T_301) begin
      ramWire_42 <= _T_298;
    end
    if (_T_308) begin
      ramWire_43 <= _T_305;
    end
    if (_T_315) begin
      ramWire_44 <= _T_312;
    end
    if (_T_322) begin
      ramWire_45 <= _T_319;
    end
    if (_T_329) begin
      ramWire_46 <= _T_326;
    end
    if (_T_336) begin
      ramWire_47 <= _T_333;
    end
    if (_T_343) begin
      ramWire_48 <= _T_340;
    end
    if (_T_350) begin
      ramWire_49 <= _T_347;
    end
    if (_T_357) begin
      ramWire_50 <= _T_354;
    end
    if (_T_364) begin
      ramWire_51 <= _T_361;
    end
    if (_T_371) begin
      ramWire_52 <= _T_368;
    end
    if (_T_378) begin
      ramWire_53 <= _T_375;
    end
    if (_T_385) begin
      ramWire_54 <= _T_382;
    end
    if (_T_392) begin
      ramWire_55 <= _T_389;
    end
    if (_T_399) begin
      ramWire_56 <= _T_396;
    end
    if (_T_406) begin
      ramWire_57 <= _T_403;
    end
    if (_T_413) begin
      ramWire_58 <= _T_410;
    end
    if (_T_420) begin
      ramWire_59 <= _T_417;
    end
    if (_T_427) begin
      ramWire_60 <= _T_424;
    end
    if (_T_434) begin
      ramWire_61 <= _T_431;
    end
    if (_T_441) begin
      ramWire_62 <= _T_438;
    end
    if (_T_448) begin
      ramWire_63 <= _T_445;
    end
  end
endmodule
module ysyx_041728(
  input         clock,
  input         reset,
  input         io_imaster_awready,
  output        io_imaster_awvalid,
  output [3:0]  io_imaster_awid,
  output [31:0] io_imaster_awaddr,
  output [7:0]  io_imaster_awlen,
  output [2:0]  io_imaster_awsize,
  output [1:0]  io_imaster_awburst,
  input         io_imaster_wready,
  output        io_imaster_wvalid,
  output [63:0] io_imaster_wdata,
  output [7:0]  io_imaster_wstrb,
  output        io_imaster_wlast,
  output        io_imaster_bready,
  input         io_imaster_bvalid,
  input  [3:0]  io_imaster_bid,
  input  [1:0]  io_imaster_bresp,
  input         io_imaster_arready,
  output        io_imaster_arvalid,
  output [3:0]  io_imaster_arid,
  output [31:0] io_imaster_araddr,
  output [7:0]  io_imaster_arlen,
  output [2:0]  io_imaster_arsize,
  output [1:0]  io_imaster_arburst,
  output        io_imaster_rready,
  input         io_imaster_rvalid,
  input  [3:0]  io_imaster_rid,
  input  [1:0]  io_imaster_rresp,
  input  [63:0] io_imaster_rdata,
  input         io_imaster_rlast,
  input         io_dmaster_awready,
  output        io_dmaster_awvalid,
  output [3:0]  io_dmaster_awid,
  output [31:0] io_dmaster_awaddr,
  output [7:0]  io_dmaster_awlen,
  output [2:0]  io_dmaster_awsize,
  output [1:0]  io_dmaster_awburst,
  input         io_dmaster_wready,
  output        io_dmaster_wvalid,
  output [63:0] io_dmaster_wdata,
  output [7:0]  io_dmaster_wstrb,
  output        io_dmaster_wlast,
  output        io_dmaster_bready,
  input         io_dmaster_bvalid,
  input  [3:0]  io_dmaster_bid,
  input  [1:0]  io_dmaster_bresp,
  input         io_dmaster_arready,
  output        io_dmaster_arvalid,
  output [3:0]  io_dmaster_arid,
  output [31:0] io_dmaster_araddr,
  output [7:0]  io_dmaster_arlen,
  output [2:0]  io_dmaster_arsize,
  output [1:0]  io_dmaster_arburst,
  output        io_dmaster_rready,
  input         io_dmaster_rvalid,
  input  [3:0]  io_dmaster_rid,
  input  [1:0]  io_dmaster_rresp,
  input  [63:0] io_dmaster_rdata,
  input         io_dmaster_rlast,
  output        io_mmio_valid,
  input         io_mmio_ready,
  input  [63:0] io_mmio_data_read,
  output [63:0] io_mmio_data_write,
  output        io_mmio_wen,
  output [31:0] io_mmio_addr,
  output [1:0]  io_mmio_rsize,
  output [7:0]  io_mmio_mask
);
  wire  riscvIns_clock; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_reset; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_io_instIO_valid; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_io_instIO_ready; // @[ysyx_22041728.scala 30:24]
  wire [63:0] riscvIns_io_instIO_data_read; // @[ysyx_22041728.scala 30:24]
  wire [31:0] riscvIns_io_instIO_addr; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_io_dataIO_valid; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_io_dataIO_ready; // @[ysyx_22041728.scala 30:24]
  wire [63:0] riscvIns_io_dataIO_data_read; // @[ysyx_22041728.scala 30:24]
  wire [63:0] riscvIns_io_dataIO_data_write; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_io_dataIO_wen; // @[ysyx_22041728.scala 30:24]
  wire [31:0] riscvIns_io_dataIO_addr; // @[ysyx_22041728.scala 30:24]
  wire [1:0] riscvIns_io_dataIO_rsize; // @[ysyx_22041728.scala 30:24]
  wire [7:0] riscvIns_io_dataIO_mask; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_intrTimeCnt_0; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_startTimeCnt; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_block2_0; // @[ysyx_22041728.scala 30:24]
  wire  riscvIns_fencei_0; // @[ysyx_22041728.scala 30:24]
  wire  iCache_clock; // @[ysyx_22041728.scala 31:22]
  wire  iCache_reset; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 31:22]
  wire [31:0] iCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 31:22]
  wire [7:0] iCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_cacheOut_r_valid_i; // @[ysyx_22041728.scala 31:22]
  wire [63:0] iCache_io_cacheOut_r_data_i; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_cacheOut_r_last_i; // @[ysyx_22041728.scala 31:22]
  wire [31:0] iCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_cacheIn_valid; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_cacheIn_ready; // @[ysyx_22041728.scala 31:22]
  wire [63:0] iCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 31:22]
  wire [31:0] iCache_io_cacheIn_addr; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 31:22]
  wire [5:0] iCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_0_rdata; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 31:22]
  wire [5:0] iCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_1_rdata; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 31:22]
  wire [5:0] iCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_2_rdata; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 31:22]
  wire  iCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 31:22]
  wire [5:0] iCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 31:22]
  wire [127:0] iCache_io_SRAMIO_3_rdata; // @[ysyx_22041728.scala 31:22]
  wire  iCache_updataICache_0; // @[ysyx_22041728.scala 31:22]
  wire  axiIIO_clock; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_reset; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_awready; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 33:22]
  wire [31:0] axiIIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 33:22]
  wire [2:0] axiIIO_io_axiIO_awsize; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_wready; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 33:22]
  wire [63:0] axiIIO_io_axiIO_wdata; // @[ysyx_22041728.scala 33:22]
  wire [7:0] axiIIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_wlast; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_bready; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_bvalid; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_arready; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 33:22]
  wire [31:0] axiIIO_io_axiIO_araddr; // @[ysyx_22041728.scala 33:22]
  wire [7:0] axiIIO_io_axiIO_arlen; // @[ysyx_22041728.scala 33:22]
  wire [2:0] axiIIO_io_axiIO_arsize; // @[ysyx_22041728.scala 33:22]
  wire [1:0] axiIIO_io_axiIO_arburst; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_rready; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_rvalid; // @[ysyx_22041728.scala 33:22]
  wire [63:0] axiIIO_io_axiIO_rdata; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_axiIO_rlast; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_cache_ar_valid_o; // @[ysyx_22041728.scala 33:22]
  wire [31:0] axiIIO_io_cache_ar_addr_o; // @[ysyx_22041728.scala 33:22]
  wire [7:0] axiIIO_io_cache_ar_len_o; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 33:22]
  wire [63:0] axiIIO_io_cache_r_data_i; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_cache_r_last_i; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_cache_w_valid_o; // @[ysyx_22041728.scala 33:22]
  wire  axiIIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 33:22]
  wire [63:0] axiIIO_io_cache_w_data_o; // @[ysyx_22041728.scala 33:22]
  wire [31:0] axiIIO_io_cache_w_addr_o; // @[ysyx_22041728.scala 33:22]
  wire [7:0] axiIIO_io_cache_w_mask_o; // @[ysyx_22041728.scala 33:22]
  wire [1:0] axiIIO_io_cache_wsize; // @[ysyx_22041728.scala 33:22]
  wire  dArbIns_io_arbIn_valid; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbIn_ready; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbIn_data_read; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbIn_data_write; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbIn_wen; // @[ysyx_22041728.scala 36:23]
  wire [31:0] dArbIns_io_arbIn_addr; // @[ysyx_22041728.scala 36:23]
  wire [1:0] dArbIns_io_arbIn_rsize; // @[ysyx_22041728.scala 36:23]
  wire [7:0] dArbIns_io_arbIn_mask; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbMMIO_valid; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbMMIO_ready; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbMMIO_data_read; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbMMIO_data_write; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbMMIO_wen; // @[ysyx_22041728.scala 36:23]
  wire [31:0] dArbIns_io_arbMMIO_addr; // @[ysyx_22041728.scala 36:23]
  wire [1:0] dArbIns_io_arbMMIO_rsize; // @[ysyx_22041728.scala 36:23]
  wire [7:0] dArbIns_io_arbMMIO_mask; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbClint_valid; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbClint_data_read; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbClint_data_write; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbClint_wen; // @[ysyx_22041728.scala 36:23]
  wire [31:0] dArbIns_io_arbClint_addr; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbDCache_valid; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbDCache_ready; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbDCache_data_read; // @[ysyx_22041728.scala 36:23]
  wire [63:0] dArbIns_io_arbDCache_data_write; // @[ysyx_22041728.scala 36:23]
  wire  dArbIns_io_arbDCache_wen; // @[ysyx_22041728.scala 36:23]
  wire [31:0] dArbIns_io_arbDCache_addr; // @[ysyx_22041728.scala 36:23]
  wire [1:0] dArbIns_io_arbDCache_rsize; // @[ysyx_22041728.scala 36:23]
  wire [7:0] dArbIns_io_arbDCache_mask; // @[ysyx_22041728.scala 36:23]
  wire  mmioDCache_clock; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_reset; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_block; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioIn_valid; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioIn_ready; // @[ysyx_22041728.scala 37:26]
  wire [63:0] mmioDCache_io_mmioIn_data_read; // @[ysyx_22041728.scala 37:26]
  wire [63:0] mmioDCache_io_mmioIn_data_write; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioIn_wen; // @[ysyx_22041728.scala 37:26]
  wire [31:0] mmioDCache_io_mmioIn_addr; // @[ysyx_22041728.scala 37:26]
  wire [1:0] mmioDCache_io_mmioIn_rsize; // @[ysyx_22041728.scala 37:26]
  wire [7:0] mmioDCache_io_mmioIn_mask; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioOut_valid; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioOut_ready; // @[ysyx_22041728.scala 37:26]
  wire [63:0] mmioDCache_io_mmioOut_data_read; // @[ysyx_22041728.scala 37:26]
  wire [63:0] mmioDCache_io_mmioOut_data_write; // @[ysyx_22041728.scala 37:26]
  wire  mmioDCache_io_mmioOut_wen; // @[ysyx_22041728.scala 37:26]
  wire [31:0] mmioDCache_io_mmioOut_addr; // @[ysyx_22041728.scala 37:26]
  wire [1:0] mmioDCache_io_mmioOut_rsize; // @[ysyx_22041728.scala 37:26]
  wire [7:0] mmioDCache_io_mmioOut_mask; // @[ysyx_22041728.scala 37:26]
  wire  dCache_clock; // @[ysyx_22041728.scala 38:22]
  wire  dCache_reset; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 38:22]
  wire [31:0] dCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 38:22]
  wire [7:0] dCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheOut_r_valid_i; // @[ysyx_22041728.scala 38:22]
  wire [63:0] dCache_io_cacheOut_r_data_i; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheOut_r_last_i; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheOut_w_valid_o; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheOut_w_ready_i; // @[ysyx_22041728.scala 38:22]
  wire [63:0] dCache_io_cacheOut_w_data_o; // @[ysyx_22041728.scala 38:22]
  wire [31:0] dCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 38:22]
  wire [7:0] dCache_io_cacheOut_w_mask_o; // @[ysyx_22041728.scala 38:22]
  wire [1:0] dCache_io_cacheOut_wsize; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheIn_valid; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheIn_ready; // @[ysyx_22041728.scala 38:22]
  wire [63:0] dCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 38:22]
  wire [63:0] dCache_io_cacheIn_data_write; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_cacheIn_wen; // @[ysyx_22041728.scala 38:22]
  wire [31:0] dCache_io_cacheIn_addr; // @[ysyx_22041728.scala 38:22]
  wire [1:0] dCache_io_cacheIn_rsize; // @[ysyx_22041728.scala 38:22]
  wire [7:0] dCache_io_cacheIn_mask; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 38:22]
  wire [5:0] dCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_0_rdata; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 38:22]
  wire [5:0] dCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_1_rdata; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 38:22]
  wire [5:0] dCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_2_rdata; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 38:22]
  wire [5:0] dCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 38:22]
  wire [127:0] dCache_io_SRAMIO_3_rdata; // @[ysyx_22041728.scala 38:22]
  wire  dCache_io_block; // @[ysyx_22041728.scala 38:22]
  wire  clintIns_clock; // @[ysyx_22041728.scala 39:25]
  wire  clintIns_reset; // @[ysyx_22041728.scala 39:25]
  wire  clintIns_io_clintIO_valid; // @[ysyx_22041728.scala 39:25]
  wire [63:0] clintIns_io_clintIO_data_read; // @[ysyx_22041728.scala 39:25]
  wire [63:0] clintIns_io_clintIO_data_write; // @[ysyx_22041728.scala 39:25]
  wire  clintIns_io_clintIO_wen; // @[ysyx_22041728.scala 39:25]
  wire [31:0] clintIns_io_clintIO_addr; // @[ysyx_22041728.scala 39:25]
  wire  clintIns_intrTimeCnt_0; // @[ysyx_22041728.scala 39:25]
  wire  clintIns_startTimeCnt_0; // @[ysyx_22041728.scala 39:25]
  wire  axiDIO_clock; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_reset; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_awready; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 45:22]
  wire [31:0] axiDIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 45:22]
  wire [2:0] axiDIO_io_axiIO_awsize; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_wready; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 45:22]
  wire [63:0] axiDIO_io_axiIO_wdata; // @[ysyx_22041728.scala 45:22]
  wire [7:0] axiDIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_wlast; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_bready; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_bvalid; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_arready; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 45:22]
  wire [31:0] axiDIO_io_axiIO_araddr; // @[ysyx_22041728.scala 45:22]
  wire [7:0] axiDIO_io_axiIO_arlen; // @[ysyx_22041728.scala 45:22]
  wire [2:0] axiDIO_io_axiIO_arsize; // @[ysyx_22041728.scala 45:22]
  wire [1:0] axiDIO_io_axiIO_arburst; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_rready; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_rvalid; // @[ysyx_22041728.scala 45:22]
  wire [63:0] axiDIO_io_axiIO_rdata; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_axiIO_rlast; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_cache_ar_valid_o; // @[ysyx_22041728.scala 45:22]
  wire [31:0] axiDIO_io_cache_ar_addr_o; // @[ysyx_22041728.scala 45:22]
  wire [7:0] axiDIO_io_cache_ar_len_o; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 45:22]
  wire [63:0] axiDIO_io_cache_r_data_i; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_cache_r_last_i; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_cache_w_valid_o; // @[ysyx_22041728.scala 45:22]
  wire  axiDIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 45:22]
  wire [63:0] axiDIO_io_cache_w_data_o; // @[ysyx_22041728.scala 45:22]
  wire [31:0] axiDIO_io_cache_w_addr_o; // @[ysyx_22041728.scala 45:22]
  wire [7:0] axiDIO_io_cache_w_mask_o; // @[ysyx_22041728.scala 45:22]
  wire [1:0] axiDIO_io_cache_wsize; // @[ysyx_22041728.scala 45:22]
  wire  mem_clock; // @[ysyx_22041728.scala 52:24]
  wire  mem_io_memIO_cen; // @[ysyx_22041728.scala 52:24]
  wire  mem_io_memIO_wen; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_io_memIO_wdata; // @[ysyx_22041728.scala 52:24]
  wire [5:0] mem_io_memIO_addr; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_io_memIO_wmask; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_io_memIO_rdata; // @[ysyx_22041728.scala 52:24]
  wire  mem_1_clock; // @[ysyx_22041728.scala 53:24]
  wire  mem_1_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  mem_1_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_1_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] mem_1_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_1_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_1_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  mem_2_clock; // @[ysyx_22041728.scala 52:24]
  wire  mem_2_io_memIO_cen; // @[ysyx_22041728.scala 52:24]
  wire  mem_2_io_memIO_wen; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_2_io_memIO_wdata; // @[ysyx_22041728.scala 52:24]
  wire [5:0] mem_2_io_memIO_addr; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_2_io_memIO_wmask; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_2_io_memIO_rdata; // @[ysyx_22041728.scala 52:24]
  wire  mem_3_clock; // @[ysyx_22041728.scala 53:24]
  wire  mem_3_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  mem_3_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_3_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] mem_3_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_3_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_3_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  mem_4_clock; // @[ysyx_22041728.scala 52:24]
  wire  mem_4_io_memIO_cen; // @[ysyx_22041728.scala 52:24]
  wire  mem_4_io_memIO_wen; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_4_io_memIO_wdata; // @[ysyx_22041728.scala 52:24]
  wire [5:0] mem_4_io_memIO_addr; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_4_io_memIO_wmask; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_4_io_memIO_rdata; // @[ysyx_22041728.scala 52:24]
  wire  mem_5_clock; // @[ysyx_22041728.scala 53:24]
  wire  mem_5_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  mem_5_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_5_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] mem_5_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_5_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_5_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  mem_6_clock; // @[ysyx_22041728.scala 52:24]
  wire  mem_6_io_memIO_cen; // @[ysyx_22041728.scala 52:24]
  wire  mem_6_io_memIO_wen; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_6_io_memIO_wdata; // @[ysyx_22041728.scala 52:24]
  wire [5:0] mem_6_io_memIO_addr; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_6_io_memIO_wmask; // @[ysyx_22041728.scala 52:24]
  wire [127:0] mem_6_io_memIO_rdata; // @[ysyx_22041728.scala 52:24]
  wire  mem_7_clock; // @[ysyx_22041728.scala 53:24]
  wire  mem_7_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  mem_7_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_7_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] mem_7_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_7_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] mem_7_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  riscv riscvIns ( // @[ysyx_22041728.scala 30:24]
    .clock(riscvIns_clock),
    .reset(riscvIns_reset),
    .io_instIO_valid(riscvIns_io_instIO_valid),
    .io_instIO_ready(riscvIns_io_instIO_ready),
    .io_instIO_data_read(riscvIns_io_instIO_data_read),
    .io_instIO_addr(riscvIns_io_instIO_addr),
    .io_dataIO_valid(riscvIns_io_dataIO_valid),
    .io_dataIO_ready(riscvIns_io_dataIO_ready),
    .io_dataIO_data_read(riscvIns_io_dataIO_data_read),
    .io_dataIO_data_write(riscvIns_io_dataIO_data_write),
    .io_dataIO_wen(riscvIns_io_dataIO_wen),
    .io_dataIO_addr(riscvIns_io_dataIO_addr),
    .io_dataIO_rsize(riscvIns_io_dataIO_rsize),
    .io_dataIO_mask(riscvIns_io_dataIO_mask),
    .intrTimeCnt_0(riscvIns_intrTimeCnt_0),
    .startTimeCnt(riscvIns_startTimeCnt),
    .block2_0(riscvIns_block2_0),
    .fencei_0(riscvIns_fencei_0)
  );
  Icache iCache ( // @[ysyx_22041728.scala 31:22]
    .clock(iCache_clock),
    .reset(iCache_reset),
    .io_cacheOut_ar_valid_o(iCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(iCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(iCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(iCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(iCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(iCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_addr_o(iCache_io_cacheOut_w_addr_o),
    .io_cacheIn_valid(iCache_io_cacheIn_valid),
    .io_cacheIn_ready(iCache_io_cacheIn_ready),
    .io_cacheIn_data_read(iCache_io_cacheIn_data_read),
    .io_cacheIn_addr(iCache_io_cacheIn_addr),
    .io_SRAMIO_0_cen(iCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(iCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(iCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(iCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(iCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(iCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(iCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(iCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(iCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(iCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(iCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(iCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(iCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(iCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(iCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(iCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(iCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(iCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(iCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(iCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(iCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(iCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(iCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(iCache_io_SRAMIO_3_rdata),
    .updataICache_0(iCache_updataICache_0)
  );
  AXICache axiIIO ( // @[ysyx_22041728.scala 33:22]
    .clock(axiIIO_clock),
    .reset(axiIIO_reset),
    .io_axiIO_awready(axiIIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiIIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiIIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiIIO_io_axiIO_awsize),
    .io_axiIO_wready(axiIIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiIIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiIIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiIIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiIIO_io_axiIO_wlast),
    .io_axiIO_bready(axiIIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiIIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiIIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiIIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiIIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiIIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiIIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiIIO_io_axiIO_arburst),
    .io_axiIO_rready(axiIIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiIIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiIIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiIIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiIIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiIIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiIIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiIIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiIIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiIIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiIIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiIIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiIIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiIIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiIIO_io_cache_w_mask_o),
    .io_cache_wsize(axiIIO_io_cache_wsize)
  );
  arbCpu2DCache dArbIns ( // @[ysyx_22041728.scala 36:23]
    .io_arbIn_valid(dArbIns_io_arbIn_valid),
    .io_arbIn_ready(dArbIns_io_arbIn_ready),
    .io_arbIn_data_read(dArbIns_io_arbIn_data_read),
    .io_arbIn_data_write(dArbIns_io_arbIn_data_write),
    .io_arbIn_wen(dArbIns_io_arbIn_wen),
    .io_arbIn_addr(dArbIns_io_arbIn_addr),
    .io_arbIn_rsize(dArbIns_io_arbIn_rsize),
    .io_arbIn_mask(dArbIns_io_arbIn_mask),
    .io_arbMMIO_valid(dArbIns_io_arbMMIO_valid),
    .io_arbMMIO_ready(dArbIns_io_arbMMIO_ready),
    .io_arbMMIO_data_read(dArbIns_io_arbMMIO_data_read),
    .io_arbMMIO_data_write(dArbIns_io_arbMMIO_data_write),
    .io_arbMMIO_wen(dArbIns_io_arbMMIO_wen),
    .io_arbMMIO_addr(dArbIns_io_arbMMIO_addr),
    .io_arbMMIO_rsize(dArbIns_io_arbMMIO_rsize),
    .io_arbMMIO_mask(dArbIns_io_arbMMIO_mask),
    .io_arbClint_valid(dArbIns_io_arbClint_valid),
    .io_arbClint_data_read(dArbIns_io_arbClint_data_read),
    .io_arbClint_data_write(dArbIns_io_arbClint_data_write),
    .io_arbClint_wen(dArbIns_io_arbClint_wen),
    .io_arbClint_addr(dArbIns_io_arbClint_addr),
    .io_arbDCache_valid(dArbIns_io_arbDCache_valid),
    .io_arbDCache_ready(dArbIns_io_arbDCache_ready),
    .io_arbDCache_data_read(dArbIns_io_arbDCache_data_read),
    .io_arbDCache_data_write(dArbIns_io_arbDCache_data_write),
    .io_arbDCache_wen(dArbIns_io_arbDCache_wen),
    .io_arbDCache_addr(dArbIns_io_arbDCache_addr),
    .io_arbDCache_rsize(dArbIns_io_arbDCache_rsize),
    .io_arbDCache_mask(dArbIns_io_arbDCache_mask)
  );
  mmioCache mmioDCache ( // @[ysyx_22041728.scala 37:26]
    .clock(mmioDCache_clock),
    .reset(mmioDCache_reset),
    .io_block(mmioDCache_io_block),
    .io_mmioIn_valid(mmioDCache_io_mmioIn_valid),
    .io_mmioIn_ready(mmioDCache_io_mmioIn_ready),
    .io_mmioIn_data_read(mmioDCache_io_mmioIn_data_read),
    .io_mmioIn_data_write(mmioDCache_io_mmioIn_data_write),
    .io_mmioIn_wen(mmioDCache_io_mmioIn_wen),
    .io_mmioIn_addr(mmioDCache_io_mmioIn_addr),
    .io_mmioIn_rsize(mmioDCache_io_mmioIn_rsize),
    .io_mmioIn_mask(mmioDCache_io_mmioIn_mask),
    .io_mmioOut_valid(mmioDCache_io_mmioOut_valid),
    .io_mmioOut_ready(mmioDCache_io_mmioOut_ready),
    .io_mmioOut_data_read(mmioDCache_io_mmioOut_data_read),
    .io_mmioOut_data_write(mmioDCache_io_mmioOut_data_write),
    .io_mmioOut_wen(mmioDCache_io_mmioOut_wen),
    .io_mmioOut_addr(mmioDCache_io_mmioOut_addr),
    .io_mmioOut_rsize(mmioDCache_io_mmioOut_rsize),
    .io_mmioOut_mask(mmioDCache_io_mmioOut_mask)
  );
  Dcache dCache ( // @[ysyx_22041728.scala 38:22]
    .clock(dCache_clock),
    .reset(dCache_reset),
    .io_cacheOut_ar_valid_o(dCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(dCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(dCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(dCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(dCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(dCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_valid_o(dCache_io_cacheOut_w_valid_o),
    .io_cacheOut_w_ready_i(dCache_io_cacheOut_w_ready_i),
    .io_cacheOut_w_data_o(dCache_io_cacheOut_w_data_o),
    .io_cacheOut_w_addr_o(dCache_io_cacheOut_w_addr_o),
    .io_cacheOut_w_mask_o(dCache_io_cacheOut_w_mask_o),
    .io_cacheOut_wsize(dCache_io_cacheOut_wsize),
    .io_cacheIn_valid(dCache_io_cacheIn_valid),
    .io_cacheIn_ready(dCache_io_cacheIn_ready),
    .io_cacheIn_data_read(dCache_io_cacheIn_data_read),
    .io_cacheIn_data_write(dCache_io_cacheIn_data_write),
    .io_cacheIn_wen(dCache_io_cacheIn_wen),
    .io_cacheIn_addr(dCache_io_cacheIn_addr),
    .io_cacheIn_rsize(dCache_io_cacheIn_rsize),
    .io_cacheIn_mask(dCache_io_cacheIn_mask),
    .io_SRAMIO_0_cen(dCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(dCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(dCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(dCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(dCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(dCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(dCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(dCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(dCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(dCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(dCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(dCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(dCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(dCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(dCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(dCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(dCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(dCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(dCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(dCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(dCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(dCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(dCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(dCache_io_SRAMIO_3_rdata),
    .io_block(dCache_io_block)
  );
  clint clintIns ( // @[ysyx_22041728.scala 39:25]
    .clock(clintIns_clock),
    .reset(clintIns_reset),
    .io_clintIO_valid(clintIns_io_clintIO_valid),
    .io_clintIO_data_read(clintIns_io_clintIO_data_read),
    .io_clintIO_data_write(clintIns_io_clintIO_data_write),
    .io_clintIO_wen(clintIns_io_clintIO_wen),
    .io_clintIO_addr(clintIns_io_clintIO_addr),
    .intrTimeCnt_0(clintIns_intrTimeCnt_0),
    .startTimeCnt_0(clintIns_startTimeCnt_0)
  );
  AXICache axiDIO ( // @[ysyx_22041728.scala 45:22]
    .clock(axiDIO_clock),
    .reset(axiDIO_reset),
    .io_axiIO_awready(axiDIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiDIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiDIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiDIO_io_axiIO_awsize),
    .io_axiIO_wready(axiDIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiDIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiDIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiDIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiDIO_io_axiIO_wlast),
    .io_axiIO_bready(axiDIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiDIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiDIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiDIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiDIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiDIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiDIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiDIO_io_axiIO_arburst),
    .io_axiIO_rready(axiDIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiDIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiDIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiDIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiDIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiDIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiDIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiDIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiDIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiDIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiDIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiDIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiDIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiDIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiDIO_io_cache_w_mask_o),
    .io_cache_wsize(axiDIO_io_cache_wsize)
  );
  mem mem ( // @[ysyx_22041728.scala 52:24]
    .clock(mem_clock),
    .io_memIO_cen(mem_io_memIO_cen),
    .io_memIO_wen(mem_io_memIO_wen),
    .io_memIO_wdata(mem_io_memIO_wdata),
    .io_memIO_addr(mem_io_memIO_addr),
    .io_memIO_wmask(mem_io_memIO_wmask),
    .io_memIO_rdata(mem_io_memIO_rdata)
  );
  mem mem_1 ( // @[ysyx_22041728.scala 53:24]
    .clock(mem_1_clock),
    .io_memIO_cen(mem_1_io_memIO_cen),
    .io_memIO_wen(mem_1_io_memIO_wen),
    .io_memIO_wdata(mem_1_io_memIO_wdata),
    .io_memIO_addr(mem_1_io_memIO_addr),
    .io_memIO_wmask(mem_1_io_memIO_wmask),
    .io_memIO_rdata(mem_1_io_memIO_rdata)
  );
  mem mem_2 ( // @[ysyx_22041728.scala 52:24]
    .clock(mem_2_clock),
    .io_memIO_cen(mem_2_io_memIO_cen),
    .io_memIO_wen(mem_2_io_memIO_wen),
    .io_memIO_wdata(mem_2_io_memIO_wdata),
    .io_memIO_addr(mem_2_io_memIO_addr),
    .io_memIO_wmask(mem_2_io_memIO_wmask),
    .io_memIO_rdata(mem_2_io_memIO_rdata)
  );
  mem mem_3 ( // @[ysyx_22041728.scala 53:24]
    .clock(mem_3_clock),
    .io_memIO_cen(mem_3_io_memIO_cen),
    .io_memIO_wen(mem_3_io_memIO_wen),
    .io_memIO_wdata(mem_3_io_memIO_wdata),
    .io_memIO_addr(mem_3_io_memIO_addr),
    .io_memIO_wmask(mem_3_io_memIO_wmask),
    .io_memIO_rdata(mem_3_io_memIO_rdata)
  );
  mem mem_4 ( // @[ysyx_22041728.scala 52:24]
    .clock(mem_4_clock),
    .io_memIO_cen(mem_4_io_memIO_cen),
    .io_memIO_wen(mem_4_io_memIO_wen),
    .io_memIO_wdata(mem_4_io_memIO_wdata),
    .io_memIO_addr(mem_4_io_memIO_addr),
    .io_memIO_wmask(mem_4_io_memIO_wmask),
    .io_memIO_rdata(mem_4_io_memIO_rdata)
  );
  mem mem_5 ( // @[ysyx_22041728.scala 53:24]
    .clock(mem_5_clock),
    .io_memIO_cen(mem_5_io_memIO_cen),
    .io_memIO_wen(mem_5_io_memIO_wen),
    .io_memIO_wdata(mem_5_io_memIO_wdata),
    .io_memIO_addr(mem_5_io_memIO_addr),
    .io_memIO_wmask(mem_5_io_memIO_wmask),
    .io_memIO_rdata(mem_5_io_memIO_rdata)
  );
  mem mem_6 ( // @[ysyx_22041728.scala 52:24]
    .clock(mem_6_clock),
    .io_memIO_cen(mem_6_io_memIO_cen),
    .io_memIO_wen(mem_6_io_memIO_wen),
    .io_memIO_wdata(mem_6_io_memIO_wdata),
    .io_memIO_addr(mem_6_io_memIO_addr),
    .io_memIO_wmask(mem_6_io_memIO_wmask),
    .io_memIO_rdata(mem_6_io_memIO_rdata)
  );
  mem mem_7 ( // @[ysyx_22041728.scala 53:24]
    .clock(mem_7_clock),
    .io_memIO_cen(mem_7_io_memIO_cen),
    .io_memIO_wen(mem_7_io_memIO_wen),
    .io_memIO_wdata(mem_7_io_memIO_wdata),
    .io_memIO_addr(mem_7_io_memIO_addr),
    .io_memIO_wmask(mem_7_io_memIO_wmask),
    .io_memIO_rdata(mem_7_io_memIO_rdata)
  );
  assign io_imaster_awvalid = axiIIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_awid = 4'h0; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_awaddr = axiIIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_awlen = 8'h0; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_awsize = axiIIO_io_axiIO_awsize; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_awburst = 2'h1; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_wvalid = axiIIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_wdata = axiIIO_io_axiIO_wdata; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_wstrb = axiIIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_wlast = axiIIO_io_axiIO_wlast; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_bready = axiIIO_io_axiIO_bready; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_arvalid = axiIIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_arid = 4'h0; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_araddr = axiIIO_io_axiIO_araddr; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_arlen = axiIIO_io_axiIO_arlen; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_arsize = axiIIO_io_axiIO_arsize; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_arburst = axiIIO_io_axiIO_arburst; // @[ysyx_22041728.scala 94:14]
  assign io_imaster_rready = axiIIO_io_axiIO_rready; // @[ysyx_22041728.scala 94:14]
  assign io_dmaster_awvalid = axiDIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_awid = 4'h0; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_awaddr = axiDIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_awlen = 8'h0; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_awsize = axiDIO_io_axiIO_awsize; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_awburst = 2'h1; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_wvalid = axiDIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_wdata = axiDIO_io_axiIO_wdata; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_wstrb = axiDIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_wlast = axiDIO_io_axiIO_wlast; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_bready = axiDIO_io_axiIO_bready; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_arvalid = axiDIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_arid = 4'h0; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_araddr = axiDIO_io_axiIO_araddr; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_arlen = axiDIO_io_axiIO_arlen; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_arsize = axiDIO_io_axiIO_arsize; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_arburst = axiDIO_io_axiIO_arburst; // @[ysyx_22041728.scala 95:14]
  assign io_dmaster_rready = axiDIO_io_axiIO_rready; // @[ysyx_22041728.scala 95:14]
  assign io_mmio_valid = mmioDCache_io_mmioOut_valid; // @[ysyx_22041728.scala 97:25]
  assign io_mmio_data_write = mmioDCache_io_mmioOut_data_write; // @[ysyx_22041728.scala 97:25]
  assign io_mmio_wen = mmioDCache_io_mmioOut_wen; // @[ysyx_22041728.scala 97:25]
  assign io_mmio_addr = mmioDCache_io_mmioOut_addr; // @[ysyx_22041728.scala 97:25]
  assign io_mmio_rsize = mmioDCache_io_mmioOut_rsize; // @[ysyx_22041728.scala 97:25]
  assign io_mmio_mask = mmioDCache_io_mmioOut_mask; // @[ysyx_22041728.scala 97:25]
  assign riscvIns_clock = clock;
  assign riscvIns_reset = reset;
  assign riscvIns_io_instIO_ready = iCache_io_cacheIn_ready; // @[ysyx_22041728.scala 32:22]
  assign riscvIns_io_instIO_data_read = iCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 32:22]
  assign riscvIns_io_dataIO_ready = dArbIns_io_arbIn_ready; // @[ysyx_22041728.scala 40:21]
  assign riscvIns_io_dataIO_data_read = dArbIns_io_arbIn_data_read; // @[ysyx_22041728.scala 40:21]
  assign riscvIns_intrTimeCnt_0 = clintIns_intrTimeCnt_0;
  assign iCache_clock = clock;
  assign iCache_reset = reset;
  assign iCache_io_cacheOut_r_valid_i = axiIIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 34:19]
  assign iCache_io_cacheOut_r_data_i = axiIIO_io_cache_r_data_i; // @[ysyx_22041728.scala 34:19]
  assign iCache_io_cacheOut_r_last_i = axiIIO_io_cache_r_last_i; // @[ysyx_22041728.scala 34:19]
  assign iCache_io_cacheIn_valid = riscvIns_io_instIO_valid; // @[ysyx_22041728.scala 32:22]
  assign iCache_io_cacheIn_addr = riscvIns_io_instIO_addr; // @[ysyx_22041728.scala 32:22]
  assign iCache_io_SRAMIO_0_rdata = mem_io_memIO_rdata; // @[ysyx_22041728.scala 54:20]
  assign iCache_io_SRAMIO_1_rdata = mem_2_io_memIO_rdata; // @[ysyx_22041728.scala 54:20]
  assign iCache_io_SRAMIO_2_rdata = mem_4_io_memIO_rdata; // @[ysyx_22041728.scala 54:20]
  assign iCache_io_SRAMIO_3_rdata = mem_6_io_memIO_rdata; // @[ysyx_22041728.scala 54:20]
  assign iCache_updataICache_0 = riscvIns_fencei_0;
  assign axiIIO_clock = clock;
  assign axiIIO_reset = reset;
  assign axiIIO_io_axiIO_awready = io_imaster_awready; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_wready = io_imaster_wready; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_bvalid = io_imaster_bvalid; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_arready = io_imaster_arready; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_rvalid = io_imaster_rvalid; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_rdata = io_imaster_rdata; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_axiIO_rlast = io_imaster_rlast; // @[ysyx_22041728.scala 94:14]
  assign axiIIO_io_cache_ar_valid_o = iCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_ar_addr_o = iCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_ar_len_o = iCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_w_valid_o = 1'h0; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_w_data_o = 64'h0; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_w_addr_o = iCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_w_mask_o = 8'h0; // @[ysyx_22041728.scala 34:19]
  assign axiIIO_io_cache_wsize = 2'h2; // @[ysyx_22041728.scala 34:19]
  assign dArbIns_io_arbIn_valid = riscvIns_io_dataIO_valid; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbIn_data_write = riscvIns_io_dataIO_data_write; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbIn_wen = riscvIns_io_dataIO_wen; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbIn_addr = riscvIns_io_dataIO_addr; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbIn_rsize = riscvIns_io_dataIO_rsize; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbIn_mask = riscvIns_io_dataIO_mask; // @[ysyx_22041728.scala 40:21]
  assign dArbIns_io_arbMMIO_ready = mmioDCache_io_mmioIn_ready; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbMMIO_data_read = mmioDCache_io_mmioIn_data_read; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbClint_data_read = clintIns_io_clintIO_data_read; // @[ysyx_22041728.scala 43:22]
  assign dArbIns_io_arbDCache_ready = dCache_io_cacheIn_ready; // @[ysyx_22041728.scala 42:24]
  assign dArbIns_io_arbDCache_data_read = dCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 42:24]
  assign mmioDCache_clock = clock;
  assign mmioDCache_reset = reset;
  assign mmioDCache_io_block = riscvIns_block2_0; // @[ysyx_22041728.scala 91:23]
  assign mmioDCache_io_mmioIn_valid = dArbIns_io_arbMMIO_valid; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioIn_data_write = dArbIns_io_arbMMIO_data_write; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioIn_wen = dArbIns_io_arbMMIO_wen; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioIn_addr = dArbIns_io_arbMMIO_addr; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioIn_rsize = dArbIns_io_arbMMIO_rsize; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioIn_mask = dArbIns_io_arbMMIO_mask; // @[ysyx_22041728.scala 41:21]
  assign mmioDCache_io_mmioOut_ready = io_mmio_ready; // @[ysyx_22041728.scala 97:25]
  assign mmioDCache_io_mmioOut_data_read = io_mmio_data_read; // @[ysyx_22041728.scala 97:25]
  assign dCache_clock = clock;
  assign dCache_reset = reset;
  assign dCache_io_cacheOut_r_valid_i = axiDIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 47:18]
  assign dCache_io_cacheOut_r_data_i = axiDIO_io_cache_r_data_i; // @[ysyx_22041728.scala 47:18]
  assign dCache_io_cacheOut_r_last_i = axiDIO_io_cache_r_last_i; // @[ysyx_22041728.scala 47:18]
  assign dCache_io_cacheOut_w_ready_i = axiDIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 47:18]
  assign dCache_io_cacheIn_valid = dArbIns_io_arbDCache_valid; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_cacheIn_data_write = dArbIns_io_arbDCache_data_write; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_cacheIn_wen = dArbIns_io_arbDCache_wen; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_cacheIn_addr = dArbIns_io_arbDCache_addr; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_cacheIn_rsize = dArbIns_io_arbDCache_rsize; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_cacheIn_mask = dArbIns_io_arbDCache_mask; // @[ysyx_22041728.scala 42:24]
  assign dCache_io_SRAMIO_0_rdata = mem_1_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign dCache_io_SRAMIO_1_rdata = mem_3_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign dCache_io_SRAMIO_2_rdata = mem_5_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign dCache_io_SRAMIO_3_rdata = mem_7_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign dCache_io_block = riscvIns_block2_0; // @[ysyx_22041728.scala 92:19]
  assign clintIns_clock = clock;
  assign clintIns_reset = reset;
  assign clintIns_io_clintIO_valid = dArbIns_io_arbClint_valid; // @[ysyx_22041728.scala 43:22]
  assign clintIns_io_clintIO_data_write = dArbIns_io_arbClint_data_write; // @[ysyx_22041728.scala 43:22]
  assign clintIns_io_clintIO_wen = dArbIns_io_arbClint_wen; // @[ysyx_22041728.scala 43:22]
  assign clintIns_io_clintIO_addr = dArbIns_io_arbClint_addr; // @[ysyx_22041728.scala 43:22]
  assign clintIns_startTimeCnt_0 = riscvIns_startTimeCnt;
  assign axiDIO_clock = clock;
  assign axiDIO_reset = reset;
  assign axiDIO_io_axiIO_awready = io_dmaster_awready; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_wready = io_dmaster_wready; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_bvalid = io_dmaster_bvalid; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_arready = io_dmaster_arready; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_rvalid = io_dmaster_rvalid; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_rdata = io_dmaster_rdata; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_axiIO_rlast = io_dmaster_rlast; // @[ysyx_22041728.scala 95:14]
  assign axiDIO_io_cache_ar_valid_o = dCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_ar_addr_o = dCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_ar_len_o = dCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_w_valid_o = dCache_io_cacheOut_w_valid_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_w_data_o = dCache_io_cacheOut_w_data_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_w_addr_o = dCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_w_mask_o = dCache_io_cacheOut_w_mask_o; // @[ysyx_22041728.scala 47:18]
  assign axiDIO_io_cache_wsize = dCache_io_cacheOut_wsize; // @[ysyx_22041728.scala 47:18]
  assign mem_clock = clock;
  assign mem_io_memIO_cen = iCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 54:20]
  assign mem_io_memIO_wen = iCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 54:20]
  assign mem_io_memIO_wdata = iCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 54:20]
  assign mem_io_memIO_addr = iCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 54:20]
  assign mem_io_memIO_wmask = iCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 54:20]
  assign mem_1_clock = clock;
  assign mem_1_io_memIO_cen = dCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 55:20]
  assign mem_1_io_memIO_wen = dCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 55:20]
  assign mem_1_io_memIO_wdata = dCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 55:20]
  assign mem_1_io_memIO_addr = dCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 55:20]
  assign mem_1_io_memIO_wmask = dCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 55:20]
  assign mem_2_clock = clock;
  assign mem_2_io_memIO_cen = iCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 54:20]
  assign mem_2_io_memIO_wen = iCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 54:20]
  assign mem_2_io_memIO_wdata = iCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 54:20]
  assign mem_2_io_memIO_addr = iCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 54:20]
  assign mem_2_io_memIO_wmask = iCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 54:20]
  assign mem_3_clock = clock;
  assign mem_3_io_memIO_cen = dCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 55:20]
  assign mem_3_io_memIO_wen = dCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 55:20]
  assign mem_3_io_memIO_wdata = dCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 55:20]
  assign mem_3_io_memIO_addr = dCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 55:20]
  assign mem_3_io_memIO_wmask = dCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 55:20]
  assign mem_4_clock = clock;
  assign mem_4_io_memIO_cen = iCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 54:20]
  assign mem_4_io_memIO_wen = iCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 54:20]
  assign mem_4_io_memIO_wdata = iCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 54:20]
  assign mem_4_io_memIO_addr = iCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 54:20]
  assign mem_4_io_memIO_wmask = iCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 54:20]
  assign mem_5_clock = clock;
  assign mem_5_io_memIO_cen = dCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 55:20]
  assign mem_5_io_memIO_wen = dCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 55:20]
  assign mem_5_io_memIO_wdata = dCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 55:20]
  assign mem_5_io_memIO_addr = dCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 55:20]
  assign mem_5_io_memIO_wmask = dCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 55:20]
  assign mem_6_clock = clock;
  assign mem_6_io_memIO_cen = iCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 54:20]
  assign mem_6_io_memIO_wen = iCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 54:20]
  assign mem_6_io_memIO_wdata = iCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 54:20]
  assign mem_6_io_memIO_addr = iCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 54:20]
  assign mem_6_io_memIO_wmask = iCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 54:20]
  assign mem_7_clock = clock;
  assign mem_7_io_memIO_cen = dCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 55:20]
  assign mem_7_io_memIO_wen = dCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 55:20]
  assign mem_7_io_memIO_wdata = dCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 55:20]
  assign mem_7_io_memIO_addr = dCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 55:20]
  assign mem_7_io_memIO_wmask = dCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 55:20]
endmodule
