module DMACtrl(
  input          clock,
  input          reset,
  input          io_dataIn_arready,
  output         io_dataIn_arvalid,
  output [31:0]  io_dataIn_araddr,
  output [7:0]   io_dataIn_arlen,
  output         io_dataIn_rready,
  input          io_dataIn_rvalid,
  input  [63:0]  io_dataIn_rdata,
  input          io_dataIn_rlast,
  output         io_dataOutMMIO_valid,
  output [63:0]  io_dataOutMMIO_data_write,
  output         io_dataOutMMIO_wen,
  output [31:0]  io_dataOutMMIO_addr,
  input          dmaEn_0,
  input  [191:0] dmaCtrl_0,
  output         blockDMA_0,
  output         DMABuzy_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] dmaSrcAddr = dmaCtrl_0[63:0]; // @[DMACtrl.scala 16:27]
  wire [63:0] dmaDstAddr = dmaCtrl_0[127:64]; // @[DMACtrl.scala 17:27]
  wire [63:0] dmaDstLen = dmaCtrl_0[191:128]; // @[DMACtrl.scala 18:26]
  reg [1:0] rState; // @[DMACtrl.scala 30:23]
  wire [1:0] idleMux = dmaEn_0 ? 2'h1 : 2'h0; // @[DMACtrl.scala 32:20]
  wire [1:0] _reqMux_T = io_dataIn_rlast ? 2'h0 : 2'h2; // @[DMACtrl.scala 35:8]
  wire  isReq = rState == 2'h1; // @[DMACtrl.scala 55:22]
  wire  isData = rState == 2'h2; // @[DMACtrl.scala 56:23]
  wire  DMABuzy = isReq | isData; // @[DMACtrl.scala 58:23]
  reg [31:0] addrCnt; // @[DMACtrl.scala 104:24]
  wire  _addrCnt_T = isData & io_dataIn_rvalid; // @[DMACtrl.scala 109:14]
  wire [31:0] _addrCnt_T_2 = addrCnt + 32'h8; // @[DMACtrl.scala 110:15]
  wire [31:0] _addrCnt_T_3 = _addrCnt_T ? _addrCnt_T_2 : addrCnt; // @[DMACtrl.scala 108:8]
  wire [63:0] _addrCnt_T_4 = isReq ? dmaDstAddr : {{32'd0}, _addrCnt_T_3}; // @[DMACtrl.scala 105:17]
  wire  blockDMA = dmaEn_0 & ~io_dataIn_rlast; // @[DMACtrl.scala 25:21]
  assign io_dataIn_arvalid = rState == 2'h1; // @[DMACtrl.scala 55:22]
  assign io_dataIn_araddr = dmaSrcAddr[31:0]; // @[DMACtrl.scala 63:20]
  assign io_dataIn_arlen = dmaDstLen[7:0]; // @[DMACtrl.scala 65:31]
  assign io_dataIn_rready = isReq | isData; // @[DMACtrl.scala 69:29]
  assign io_dataOutMMIO_valid = DMABuzy & io_dataIn_rvalid; // @[DMACtrl.scala 71:45]
  assign io_dataOutMMIO_data_write = io_dataIn_rdata; // @[DMACtrl.scala 73:29]
  assign io_dataOutMMIO_wen = isData & io_dataIn_rvalid; // @[DMACtrl.scala 116:32]
  assign io_dataOutMMIO_addr = addrCnt; // @[DMACtrl.scala 114:23]
  assign blockDMA_0 = blockDMA;
  assign DMABuzy_0 = DMABuzy;
  always @(posedge clock) begin
    if (reset) begin // @[DMACtrl.scala 30:23]
      rState <= 2'h0; // @[DMACtrl.scala 30:23]
    end else if (2'h2 == rState) begin // @[Mux.scala 80:57]
      rState <= _reqMux_T;
    end else if (2'h1 == rState) begin // @[Mux.scala 80:57]
      if (io_dataIn_arready) begin // @[DMACtrl.scala 33:19]
        rState <= _reqMux_T;
      end else begin
        rState <= 2'h1;
      end
    end else if (2'h0 == rState) begin // @[Mux.scala 80:57]
      rState <= idleMux;
    end
    if (reset) begin // @[DMACtrl.scala 104:24]
      addrCnt <= 32'h0; // @[DMACtrl.scala 104:24]
    end else begin
      addrCnt <= _addrCnt_T_4[31:0]; // @[DMACtrl.scala 105:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  addrCnt = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module iFetch(
  input         clock,
  input         reset,
  input  [31:0] io_instIn,
  output [31:0] io_instOut,
  output [31:0] io_pc,
  output [31:0] io_snpc,
  input  [31:0] io_dnpc,
  input         io_jump,
  input         intrTimeCnt_0,
  input         hazardPCBlock_0,
  input         blockDMA_0,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[Reg.scala 27:20]
  wire [31:0] snpc = pc + 32'h4; // @[iFetch.scala 40:14]
  wire  _pc_T_6 = ~(block1_0 | block23_0 | blockDMA_0) & (~hazardPCBlock_0 | intrTimeCnt_0); // @[iFetch.scala 38:101]
  assign io_instOut = io_instIn; // @[iFetch.scala 55:14]
  assign io_pc = pc; // @[iFetch.scala 48:9]
  assign io_snpc = pc + 32'h4; // @[iFetch.scala 40:14]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      pc <= 32'h80000000; // @[Reg.scala 27:20]
    end else if (_pc_T_6) begin // @[Reg.scala 28:19]
      if (io_jump) begin // @[iFetch.scala 38:25]
        pc <= io_dnpc;
      end else begin
        pc <= snpc;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module immeGen(
  input  [31:0] io_inst,
  output [63:0] io_imme
);
  wire [11:0] Iimm_lo = io_inst[31:20]; // @[immeGen.scala 40:31]
  wire  Iimm_signBit = Iimm_lo[11]; // @[immeGen.scala 17:22]
  wire [51:0] Iimm_hi = Iimm_signBit ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Iimm = {Iimm_hi,Iimm_lo}; // @[Cat.scala 30:58]
  wire [6:0] Simm_hi = io_inst[31:25]; // @[immeGen.scala 41:35]
  wire [4:0] Simm_lo = io_inst[11:7]; // @[immeGen.scala 41:52]
  wire [11:0] Simm_lo_1 = {Simm_hi,Simm_lo}; // @[Cat.scala 30:58]
  wire  Simm_signBit = Simm_lo_1[11]; // @[immeGen.scala 17:22]
  wire [51:0] Simm_hi_1 = Simm_signBit ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Simm = {Simm_hi_1,Simm_hi,Simm_lo}; // @[Cat.scala 30:58]
  wire  Bimm_hi_hi_hi = io_inst[31]; // @[immeGen.scala 42:35]
  wire  Bimm_hi_hi_lo = io_inst[7]; // @[immeGen.scala 42:48]
  wire [5:0] Bimm_hi_lo = io_inst[30:25]; // @[immeGen.scala 42:60]
  wire [3:0] Bimm_lo_hi = io_inst[11:8]; // @[immeGen.scala 42:77]
  wire [12:0] Bimm_lo_1 = {Bimm_hi_hi_hi,Bimm_hi_hi_lo,Bimm_hi_lo,Bimm_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  Bimm_signBit = Bimm_lo_1[12]; // @[immeGen.scala 17:22]
  wire [50:0] Bimm_hi_1 = Bimm_signBit ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Bimm = {Bimm_hi_1,Bimm_hi_hi_hi,Bimm_hi_hi_lo,Bimm_hi_lo,Bimm_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] Uimm_hi = io_inst[31:12]; // @[immeGen.scala 43:35]
  wire [31:0] Uimm_lo = {Uimm_hi,12'h0}; // @[Cat.scala 30:58]
  wire  Uimm_signBit = Uimm_lo[31]; // @[immeGen.scala 17:22]
  wire [31:0] Uimm_hi_1 = Uimm_signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Uimm = {Uimm_hi_1,Uimm_hi,12'h0}; // @[Cat.scala 30:58]
  wire [7:0] Jimm_hi_hi_lo = io_inst[19:12]; // @[immeGen.scala 44:48]
  wire  Jimm_hi_lo = io_inst[20]; // @[immeGen.scala 44:65]
  wire [9:0] Jimm_lo_hi = io_inst[30:21]; // @[immeGen.scala 44:78]
  wire [20:0] Jimm_lo_1 = {Bimm_hi_hi_hi,Jimm_hi_hi_lo,Jimm_hi_lo,Jimm_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire  Jimm_signBit = Jimm_lo_1[20]; // @[immeGen.scala 17:22]
  wire [42:0] Jimm_hi_1 = Jimm_signBit ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] Jimm = {Jimm_hi_1,Bimm_hi_hi_hi,Jimm_hi_hi_lo,Jimm_hi_lo,Jimm_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T = io_inst & 32'hfc00707f; // @[immeGen.scala 51:47]
  wire  _T_1 = 32'h1013 == _T; // @[immeGen.scala 51:47]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[immeGen.scala 51:47]
  wire  _T_3 = 32'h13 == _T_2; // @[immeGen.scala 51:47]
  wire [31:0] _T_4 = io_inst & 32'hfe00707f; // @[immeGen.scala 51:47]
  wire  _T_5 = 32'h101b == _T_4; // @[immeGen.scala 51:47]
  wire  _T_7 = 32'h5013 == _T; // @[immeGen.scala 51:47]
  wire  _T_9 = 32'h6063 == _T_2; // @[immeGen.scala 55:47]
  wire  _T_11 = 32'h6013 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_13 = 32'h7013 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_15 = 32'h4063 == _T_2; // @[immeGen.scala 55:47]
  wire  _T_17 = 32'h501b == _T_4; // @[immeGen.scala 51:47]
  wire  _T_19 = 32'h3003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_21 = 32'h3013 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_23 = 32'h1003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_25 = 32'h4000501b == _T_4; // @[immeGen.scala 51:47]
  wire  _T_27 = 32'h67 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_29 = 32'h1063 == _T_2; // @[immeGen.scala 55:47]
  wire  _T_31 = 32'h1b == _T_2; // @[immeGen.scala 51:47]
  wire  _T_33 = 32'h3023 == _T_2; // @[immeGen.scala 54:47]
  wire  _T_35 = 32'h4013 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_37 = 32'h2003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_39 = 32'h4003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_41 = 32'h5003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_43 = 32'h3 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_45 = 32'h7063 == _T_2; // @[immeGen.scala 55:47]
  wire  _T_47 = 32'h23 == _T_2; // @[immeGen.scala 54:47]
  wire  _T_49 = 32'h2023 == _T_2; // @[immeGen.scala 54:47]
  wire  _T_51 = 32'h40005013 == _T; // @[immeGen.scala 51:47]
  wire  _T_53 = 32'h63 == _T_2; // @[immeGen.scala 55:47]
  wire  _T_55 = 32'h5063 == _T_2; // @[immeGen.scala 55:47]
  wire [31:0] _T_56 = io_inst & 32'h7f; // @[immeGen.scala 53:47]
  wire  _T_57 = 32'h17 == _T_56; // @[immeGen.scala 53:47]
  wire  _T_59 = 32'h6003 == _T_2; // @[immeGen.scala 51:47]
  wire  _T_61 = 32'h37 == _T_56; // @[immeGen.scala 53:47]
  wire  _T_63 = 32'h1023 == _T_2; // @[immeGen.scala 54:47]
  wire  _T_65 = 32'h6f == _T_56; // @[immeGen.scala 52:47]
  wire  _T_67 = 32'h1073 == _T_2; // @[immeGen.scala 61:29]
  wire  _T_69 = 32'h2073 == _T_2; // @[immeGen.scala 62:29]
  wire  _T_71 = 32'h6073 == _T_2; // @[immeGen.scala 63:29]
  wire  _T_73 = 32'h7073 == _T_2; // @[immeGen.scala 64:29]
  wire  _T_75 = 32'h3073 == _T_2; // @[immeGen.scala 65:29]
  wire [63:0] _io_imme_T = _T_75 ? Iimm : 64'h0; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_1 = _T_73 ? Iimm : _io_imme_T; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_2 = _T_71 ? Iimm : _io_imme_T_1; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_3 = _T_69 ? Iimm : _io_imme_T_2; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_4 = _T_67 ? Iimm : _io_imme_T_3; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_5 = _T_65 ? Jimm : _io_imme_T_4; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_6 = _T_63 ? Simm : _io_imme_T_5; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_7 = _T_61 ? Uimm : _io_imme_T_6; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_8 = _T_59 ? Iimm : _io_imme_T_7; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_9 = _T_57 ? Uimm : _io_imme_T_8; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_10 = _T_55 ? Bimm : _io_imme_T_9; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_11 = _T_53 ? Bimm : _io_imme_T_10; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_12 = _T_51 ? Iimm : _io_imme_T_11; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_13 = _T_49 ? Simm : _io_imme_T_12; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_14 = _T_47 ? Simm : _io_imme_T_13; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_15 = _T_45 ? Bimm : _io_imme_T_14; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_16 = _T_43 ? Iimm : _io_imme_T_15; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_17 = _T_41 ? Iimm : _io_imme_T_16; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_18 = _T_39 ? Iimm : _io_imme_T_17; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_19 = _T_37 ? Iimm : _io_imme_T_18; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_20 = _T_35 ? Iimm : _io_imme_T_19; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_21 = _T_33 ? Simm : _io_imme_T_20; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_22 = _T_31 ? Iimm : _io_imme_T_21; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_23 = _T_29 ? Bimm : _io_imme_T_22; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_24 = _T_27 ? Iimm : _io_imme_T_23; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_25 = _T_25 ? Iimm : _io_imme_T_24; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_26 = _T_23 ? Iimm : _io_imme_T_25; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_27 = _T_21 ? Iimm : _io_imme_T_26; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_28 = _T_19 ? Iimm : _io_imme_T_27; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_29 = _T_17 ? Iimm : _io_imme_T_28; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_30 = _T_15 ? Bimm : _io_imme_T_29; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_31 = _T_13 ? Iimm : _io_imme_T_30; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_32 = _T_11 ? Iimm : _io_imme_T_31; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_33 = _T_9 ? Bimm : _io_imme_T_32; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_34 = _T_7 ? Iimm : _io_imme_T_33; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_35 = _T_5 ? Iimm : _io_imme_T_34; // @[Mux.scala 98:16]
  wire [63:0] _io_imme_T_36 = _T_3 ? Iimm : _io_imme_T_35; // @[Mux.scala 98:16]
  assign io_imme = _T_1 ? Iimm : _io_imme_T_36; // @[Mux.scala 98:16]
endmodule
module RF(
  input         clock,
  input  [31:0] io_pc,
  input         io_we,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_rd,
  input  [4:0]  io_rdID,
  output [63:0] io_dout1,
  output [63:0] io_dout2,
  output [63:0] io_rdDout,
  input  [63:0] io_din,
  input  [4:0]  io_rsWB,
  output [63:0] io_doutWB,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] DPIC_RegRead_ins_inst_0; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_1; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_2; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_3; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_4; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_5; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_6; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_7; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_8; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_9; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_10; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_11; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_12; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_13; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_14; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_15; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_16; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_17; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_18; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_19; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_20; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_21; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_22; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_23; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_24; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_25; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_26; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_27; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_28; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_29; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_30; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_inst_31; // @[regFile.scala 29:32]
  wire [63:0] DPIC_RegRead_ins_pc; // @[regFile.scala 29:32]
  wire  en = io_we & io_rd == 5'h1; // @[regFile.scala 54:13]
  wire  _regData_T_7 = en & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_1; // @[Reg.scala 15:16]
  wire  en_1 = io_we & io_rd == 5'h2; // @[regFile.scala 54:13]
  wire  _regData_T_11 = en_1 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_2; // @[Reg.scala 15:16]
  wire  en_2 = io_we & io_rd == 5'h3; // @[regFile.scala 54:13]
  wire  _regData_T_15 = en_2 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_3; // @[Reg.scala 15:16]
  wire  en_3 = io_we & io_rd == 5'h4; // @[regFile.scala 54:13]
  wire  _regData_T_19 = en_3 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_4; // @[Reg.scala 15:16]
  wire  en_4 = io_we & io_rd == 5'h5; // @[regFile.scala 54:13]
  wire  _regData_T_23 = en_4 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_5; // @[Reg.scala 15:16]
  wire  en_5 = io_we & io_rd == 5'h6; // @[regFile.scala 54:13]
  wire  _regData_T_27 = en_5 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_6; // @[Reg.scala 15:16]
  wire  en_6 = io_we & io_rd == 5'h7; // @[regFile.scala 54:13]
  wire  _regData_T_31 = en_6 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_7; // @[Reg.scala 15:16]
  wire  en_7 = io_we & io_rd == 5'h8; // @[regFile.scala 54:13]
  wire  _regData_T_35 = en_7 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_8; // @[Reg.scala 15:16]
  wire  en_8 = io_we & io_rd == 5'h9; // @[regFile.scala 54:13]
  wire  _regData_T_39 = en_8 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_9; // @[Reg.scala 15:16]
  wire  en_9 = io_we & io_rd == 5'ha; // @[regFile.scala 54:13]
  wire  _regData_T_43 = en_9 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_10; // @[Reg.scala 15:16]
  wire  en_10 = io_we & io_rd == 5'hb; // @[regFile.scala 54:13]
  wire  _regData_T_47 = en_10 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_11; // @[Reg.scala 15:16]
  wire  en_11 = io_we & io_rd == 5'hc; // @[regFile.scala 54:13]
  wire  _regData_T_51 = en_11 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_12; // @[Reg.scala 15:16]
  wire  en_12 = io_we & io_rd == 5'hd; // @[regFile.scala 54:13]
  wire  _regData_T_55 = en_12 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_13; // @[Reg.scala 15:16]
  wire  en_13 = io_we & io_rd == 5'he; // @[regFile.scala 54:13]
  wire  _regData_T_59 = en_13 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_14; // @[Reg.scala 15:16]
  wire  en_14 = io_we & io_rd == 5'hf; // @[regFile.scala 54:13]
  wire  _regData_T_63 = en_14 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_15; // @[Reg.scala 15:16]
  wire  en_15 = io_we & io_rd == 5'h10; // @[regFile.scala 54:13]
  wire  _regData_T_67 = en_15 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_16; // @[Reg.scala 15:16]
  wire  en_16 = io_we & io_rd == 5'h11; // @[regFile.scala 54:13]
  wire  _regData_T_71 = en_16 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_17; // @[Reg.scala 15:16]
  wire  en_17 = io_we & io_rd == 5'h12; // @[regFile.scala 54:13]
  wire  _regData_T_75 = en_17 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_18; // @[Reg.scala 15:16]
  wire  en_18 = io_we & io_rd == 5'h13; // @[regFile.scala 54:13]
  wire  _regData_T_79 = en_18 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_19; // @[Reg.scala 15:16]
  wire  en_19 = io_we & io_rd == 5'h14; // @[regFile.scala 54:13]
  wire  _regData_T_83 = en_19 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_20; // @[Reg.scala 15:16]
  wire  en_20 = io_we & io_rd == 5'h15; // @[regFile.scala 54:13]
  wire  _regData_T_87 = en_20 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_21; // @[Reg.scala 15:16]
  wire  en_21 = io_we & io_rd == 5'h16; // @[regFile.scala 54:13]
  wire  _regData_T_91 = en_21 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_22; // @[Reg.scala 15:16]
  wire  en_22 = io_we & io_rd == 5'h17; // @[regFile.scala 54:13]
  wire  _regData_T_95 = en_22 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_23; // @[Reg.scala 15:16]
  wire  en_23 = io_we & io_rd == 5'h18; // @[regFile.scala 54:13]
  wire  _regData_T_99 = en_23 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_24; // @[Reg.scala 15:16]
  wire  en_24 = io_we & io_rd == 5'h19; // @[regFile.scala 54:13]
  wire  _regData_T_103 = en_24 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_25; // @[Reg.scala 15:16]
  wire  en_25 = io_we & io_rd == 5'h1a; // @[regFile.scala 54:13]
  wire  _regData_T_107 = en_25 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_26; // @[Reg.scala 15:16]
  wire  en_26 = io_we & io_rd == 5'h1b; // @[regFile.scala 54:13]
  wire  _regData_T_111 = en_26 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_27; // @[Reg.scala 15:16]
  wire  en_27 = io_we & io_rd == 5'h1c; // @[regFile.scala 54:13]
  wire  _regData_T_115 = en_27 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_28; // @[Reg.scala 15:16]
  wire  en_28 = io_we & io_rd == 5'h1d; // @[regFile.scala 54:13]
  wire  _regData_T_119 = en_28 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_29; // @[Reg.scala 15:16]
  wire  en_29 = io_we & io_rd == 5'h1e; // @[regFile.scala 54:13]
  wire  _regData_T_123 = en_29 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_30; // @[Reg.scala 15:16]
  wire  en_30 = io_we & io_rd == 5'h1f; // @[regFile.scala 54:13]
  wire  _regData_T_127 = en_30 & ~(block1_0 | block23_0 | block23_0); // @[regFile.scala 66:38]
  reg [63:0] regData_r_31; // @[Reg.scala 15:16]
  wire [63:0] _io_dout1_T_1 = 5'h1 == io_rs1 ? regData_r_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_3 = 5'h2 == io_rs1 ? regData_r_2 : _io_dout1_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_5 = 5'h3 == io_rs1 ? regData_r_3 : _io_dout1_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_7 = 5'h4 == io_rs1 ? regData_r_4 : _io_dout1_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_9 = 5'h5 == io_rs1 ? regData_r_5 : _io_dout1_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_11 = 5'h6 == io_rs1 ? regData_r_6 : _io_dout1_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_13 = 5'h7 == io_rs1 ? regData_r_7 : _io_dout1_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_15 = 5'h8 == io_rs1 ? regData_r_8 : _io_dout1_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_17 = 5'h9 == io_rs1 ? regData_r_9 : _io_dout1_T_15; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_19 = 5'ha == io_rs1 ? regData_r_10 : _io_dout1_T_17; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_21 = 5'hb == io_rs1 ? regData_r_11 : _io_dout1_T_19; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_23 = 5'hc == io_rs1 ? regData_r_12 : _io_dout1_T_21; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_25 = 5'hd == io_rs1 ? regData_r_13 : _io_dout1_T_23; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_27 = 5'he == io_rs1 ? regData_r_14 : _io_dout1_T_25; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_29 = 5'hf == io_rs1 ? regData_r_15 : _io_dout1_T_27; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_31 = 5'h10 == io_rs1 ? regData_r_16 : _io_dout1_T_29; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_33 = 5'h11 == io_rs1 ? regData_r_17 : _io_dout1_T_31; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_35 = 5'h12 == io_rs1 ? regData_r_18 : _io_dout1_T_33; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_37 = 5'h13 == io_rs1 ? regData_r_19 : _io_dout1_T_35; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_39 = 5'h14 == io_rs1 ? regData_r_20 : _io_dout1_T_37; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_41 = 5'h15 == io_rs1 ? regData_r_21 : _io_dout1_T_39; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_43 = 5'h16 == io_rs1 ? regData_r_22 : _io_dout1_T_41; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_45 = 5'h17 == io_rs1 ? regData_r_23 : _io_dout1_T_43; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_47 = 5'h18 == io_rs1 ? regData_r_24 : _io_dout1_T_45; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_49 = 5'h19 == io_rs1 ? regData_r_25 : _io_dout1_T_47; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_51 = 5'h1a == io_rs1 ? regData_r_26 : _io_dout1_T_49; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_53 = 5'h1b == io_rs1 ? regData_r_27 : _io_dout1_T_51; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_55 = 5'h1c == io_rs1 ? regData_r_28 : _io_dout1_T_53; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_57 = 5'h1d == io_rs1 ? regData_r_29 : _io_dout1_T_55; // @[Mux.scala 80:57]
  wire [63:0] _io_dout1_T_59 = 5'h1e == io_rs1 ? regData_r_30 : _io_dout1_T_57; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_1 = 5'h1 == io_rs2 ? regData_r_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_3 = 5'h2 == io_rs2 ? regData_r_2 : _io_dout2_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_5 = 5'h3 == io_rs2 ? regData_r_3 : _io_dout2_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_7 = 5'h4 == io_rs2 ? regData_r_4 : _io_dout2_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_9 = 5'h5 == io_rs2 ? regData_r_5 : _io_dout2_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_11 = 5'h6 == io_rs2 ? regData_r_6 : _io_dout2_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_13 = 5'h7 == io_rs2 ? regData_r_7 : _io_dout2_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_15 = 5'h8 == io_rs2 ? regData_r_8 : _io_dout2_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_17 = 5'h9 == io_rs2 ? regData_r_9 : _io_dout2_T_15; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_19 = 5'ha == io_rs2 ? regData_r_10 : _io_dout2_T_17; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_21 = 5'hb == io_rs2 ? regData_r_11 : _io_dout2_T_19; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_23 = 5'hc == io_rs2 ? regData_r_12 : _io_dout2_T_21; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_25 = 5'hd == io_rs2 ? regData_r_13 : _io_dout2_T_23; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_27 = 5'he == io_rs2 ? regData_r_14 : _io_dout2_T_25; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_29 = 5'hf == io_rs2 ? regData_r_15 : _io_dout2_T_27; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_31 = 5'h10 == io_rs2 ? regData_r_16 : _io_dout2_T_29; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_33 = 5'h11 == io_rs2 ? regData_r_17 : _io_dout2_T_31; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_35 = 5'h12 == io_rs2 ? regData_r_18 : _io_dout2_T_33; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_37 = 5'h13 == io_rs2 ? regData_r_19 : _io_dout2_T_35; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_39 = 5'h14 == io_rs2 ? regData_r_20 : _io_dout2_T_37; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_41 = 5'h15 == io_rs2 ? regData_r_21 : _io_dout2_T_39; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_43 = 5'h16 == io_rs2 ? regData_r_22 : _io_dout2_T_41; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_45 = 5'h17 == io_rs2 ? regData_r_23 : _io_dout2_T_43; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_47 = 5'h18 == io_rs2 ? regData_r_24 : _io_dout2_T_45; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_49 = 5'h19 == io_rs2 ? regData_r_25 : _io_dout2_T_47; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_51 = 5'h1a == io_rs2 ? regData_r_26 : _io_dout2_T_49; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_53 = 5'h1b == io_rs2 ? regData_r_27 : _io_dout2_T_51; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_55 = 5'h1c == io_rs2 ? regData_r_28 : _io_dout2_T_53; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_57 = 5'h1d == io_rs2 ? regData_r_29 : _io_dout2_T_55; // @[Mux.scala 80:57]
  wire [63:0] _io_dout2_T_59 = 5'h1e == io_rs2 ? regData_r_30 : _io_dout2_T_57; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_1 = 5'h1 == io_rdID ? regData_r_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_3 = 5'h2 == io_rdID ? regData_r_2 : _io_rdDout_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_5 = 5'h3 == io_rdID ? regData_r_3 : _io_rdDout_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_7 = 5'h4 == io_rdID ? regData_r_4 : _io_rdDout_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_9 = 5'h5 == io_rdID ? regData_r_5 : _io_rdDout_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_11 = 5'h6 == io_rdID ? regData_r_6 : _io_rdDout_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_13 = 5'h7 == io_rdID ? regData_r_7 : _io_rdDout_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_15 = 5'h8 == io_rdID ? regData_r_8 : _io_rdDout_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_17 = 5'h9 == io_rdID ? regData_r_9 : _io_rdDout_T_15; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_19 = 5'ha == io_rdID ? regData_r_10 : _io_rdDout_T_17; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_21 = 5'hb == io_rdID ? regData_r_11 : _io_rdDout_T_19; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_23 = 5'hc == io_rdID ? regData_r_12 : _io_rdDout_T_21; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_25 = 5'hd == io_rdID ? regData_r_13 : _io_rdDout_T_23; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_27 = 5'he == io_rdID ? regData_r_14 : _io_rdDout_T_25; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_29 = 5'hf == io_rdID ? regData_r_15 : _io_rdDout_T_27; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_31 = 5'h10 == io_rdID ? regData_r_16 : _io_rdDout_T_29; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_33 = 5'h11 == io_rdID ? regData_r_17 : _io_rdDout_T_31; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_35 = 5'h12 == io_rdID ? regData_r_18 : _io_rdDout_T_33; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_37 = 5'h13 == io_rdID ? regData_r_19 : _io_rdDout_T_35; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_39 = 5'h14 == io_rdID ? regData_r_20 : _io_rdDout_T_37; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_41 = 5'h15 == io_rdID ? regData_r_21 : _io_rdDout_T_39; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_43 = 5'h16 == io_rdID ? regData_r_22 : _io_rdDout_T_41; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_45 = 5'h17 == io_rdID ? regData_r_23 : _io_rdDout_T_43; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_47 = 5'h18 == io_rdID ? regData_r_24 : _io_rdDout_T_45; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_49 = 5'h19 == io_rdID ? regData_r_25 : _io_rdDout_T_47; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_51 = 5'h1a == io_rdID ? regData_r_26 : _io_rdDout_T_49; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_53 = 5'h1b == io_rdID ? regData_r_27 : _io_rdDout_T_51; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_55 = 5'h1c == io_rdID ? regData_r_28 : _io_rdDout_T_53; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_57 = 5'h1d == io_rdID ? regData_r_29 : _io_rdDout_T_55; // @[Mux.scala 80:57]
  wire [63:0] _io_rdDout_T_59 = 5'h1e == io_rdID ? regData_r_30 : _io_rdDout_T_57; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_1 = 5'h1 == io_rsWB ? regData_r_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_3 = 5'h2 == io_rsWB ? regData_r_2 : _io_doutWB_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_5 = 5'h3 == io_rsWB ? regData_r_3 : _io_doutWB_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_7 = 5'h4 == io_rsWB ? regData_r_4 : _io_doutWB_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_9 = 5'h5 == io_rsWB ? regData_r_5 : _io_doutWB_T_7; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_11 = 5'h6 == io_rsWB ? regData_r_6 : _io_doutWB_T_9; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_13 = 5'h7 == io_rsWB ? regData_r_7 : _io_doutWB_T_11; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_15 = 5'h8 == io_rsWB ? regData_r_8 : _io_doutWB_T_13; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_17 = 5'h9 == io_rsWB ? regData_r_9 : _io_doutWB_T_15; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_19 = 5'ha == io_rsWB ? regData_r_10 : _io_doutWB_T_17; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_21 = 5'hb == io_rsWB ? regData_r_11 : _io_doutWB_T_19; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_23 = 5'hc == io_rsWB ? regData_r_12 : _io_doutWB_T_21; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_25 = 5'hd == io_rsWB ? regData_r_13 : _io_doutWB_T_23; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_27 = 5'he == io_rsWB ? regData_r_14 : _io_doutWB_T_25; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_29 = 5'hf == io_rsWB ? regData_r_15 : _io_doutWB_T_27; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_31 = 5'h10 == io_rsWB ? regData_r_16 : _io_doutWB_T_29; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_33 = 5'h11 == io_rsWB ? regData_r_17 : _io_doutWB_T_31; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_35 = 5'h12 == io_rsWB ? regData_r_18 : _io_doutWB_T_33; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_37 = 5'h13 == io_rsWB ? regData_r_19 : _io_doutWB_T_35; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_39 = 5'h14 == io_rsWB ? regData_r_20 : _io_doutWB_T_37; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_41 = 5'h15 == io_rsWB ? regData_r_21 : _io_doutWB_T_39; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_43 = 5'h16 == io_rsWB ? regData_r_22 : _io_doutWB_T_41; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_45 = 5'h17 == io_rsWB ? regData_r_23 : _io_doutWB_T_43; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_47 = 5'h18 == io_rsWB ? regData_r_24 : _io_doutWB_T_45; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_49 = 5'h19 == io_rsWB ? regData_r_25 : _io_doutWB_T_47; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_51 = 5'h1a == io_rsWB ? regData_r_26 : _io_doutWB_T_49; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_53 = 5'h1b == io_rsWB ? regData_r_27 : _io_doutWB_T_51; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_55 = 5'h1c == io_rsWB ? regData_r_28 : _io_doutWB_T_53; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_57 = 5'h1d == io_rsWB ? regData_r_29 : _io_doutWB_T_55; // @[Mux.scala 80:57]
  wire [63:0] _io_doutWB_T_59 = 5'h1e == io_rsWB ? regData_r_30 : _io_doutWB_T_57; // @[Mux.scala 80:57]
  DPIC_RegRead DPIC_RegRead_ins ( // @[regFile.scala 29:32]
    .inst_0(DPIC_RegRead_ins_inst_0),
    .inst_1(DPIC_RegRead_ins_inst_1),
    .inst_2(DPIC_RegRead_ins_inst_2),
    .inst_3(DPIC_RegRead_ins_inst_3),
    .inst_4(DPIC_RegRead_ins_inst_4),
    .inst_5(DPIC_RegRead_ins_inst_5),
    .inst_6(DPIC_RegRead_ins_inst_6),
    .inst_7(DPIC_RegRead_ins_inst_7),
    .inst_8(DPIC_RegRead_ins_inst_8),
    .inst_9(DPIC_RegRead_ins_inst_9),
    .inst_10(DPIC_RegRead_ins_inst_10),
    .inst_11(DPIC_RegRead_ins_inst_11),
    .inst_12(DPIC_RegRead_ins_inst_12),
    .inst_13(DPIC_RegRead_ins_inst_13),
    .inst_14(DPIC_RegRead_ins_inst_14),
    .inst_15(DPIC_RegRead_ins_inst_15),
    .inst_16(DPIC_RegRead_ins_inst_16),
    .inst_17(DPIC_RegRead_ins_inst_17),
    .inst_18(DPIC_RegRead_ins_inst_18),
    .inst_19(DPIC_RegRead_ins_inst_19),
    .inst_20(DPIC_RegRead_ins_inst_20),
    .inst_21(DPIC_RegRead_ins_inst_21),
    .inst_22(DPIC_RegRead_ins_inst_22),
    .inst_23(DPIC_RegRead_ins_inst_23),
    .inst_24(DPIC_RegRead_ins_inst_24),
    .inst_25(DPIC_RegRead_ins_inst_25),
    .inst_26(DPIC_RegRead_ins_inst_26),
    .inst_27(DPIC_RegRead_ins_inst_27),
    .inst_28(DPIC_RegRead_ins_inst_28),
    .inst_29(DPIC_RegRead_ins_inst_29),
    .inst_30(DPIC_RegRead_ins_inst_30),
    .inst_31(DPIC_RegRead_ins_inst_31),
    .pc(DPIC_RegRead_ins_pc)
  );
  assign io_dout1 = 5'h1f == io_rs1 ? regData_r_31 : _io_dout1_T_59; // @[Mux.scala 80:57]
  assign io_dout2 = 5'h1f == io_rs2 ? regData_r_31 : _io_dout2_T_59; // @[Mux.scala 80:57]
  assign io_rdDout = 5'h1f == io_rdID ? regData_r_31 : _io_rdDout_T_59; // @[Mux.scala 80:57]
  assign io_doutWB = 5'h1f == io_rsWB ? regData_r_31 : _io_doutWB_T_59; // @[Mux.scala 80:57]
  assign DPIC_RegRead_ins_inst_0 = 64'h0; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_1 = regData_r_1; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_2 = regData_r_2; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_3 = regData_r_3; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_4 = regData_r_4; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_5 = regData_r_5; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_6 = regData_r_6; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_7 = regData_r_7; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_8 = regData_r_8; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_9 = regData_r_9; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_10 = regData_r_10; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_11 = regData_r_11; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_12 = regData_r_12; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_13 = regData_r_13; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_14 = regData_r_14; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_15 = regData_r_15; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_16 = regData_r_16; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_17 = regData_r_17; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_18 = regData_r_18; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_19 = regData_r_19; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_20 = regData_r_20; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_21 = regData_r_21; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_22 = regData_r_22; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_23 = regData_r_23; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_24 = regData_r_24; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_25 = regData_r_25; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_26 = regData_r_26; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_27 = regData_r_27; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_28 = regData_r_28; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_29 = regData_r_29; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_30 = regData_r_30; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_inst_31 = regData_r_31; // @[regFile.scala 50:23 regFile.scala 66:13]
  assign DPIC_RegRead_ins_pc = {{32'd0}, io_pc}; // @[regFile.scala 30:26]
  always @(posedge clock) begin
    if (_regData_T_7) begin // @[Reg.scala 16:19]
      regData_r_1 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_11) begin // @[Reg.scala 16:19]
      regData_r_2 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_15) begin // @[Reg.scala 16:19]
      regData_r_3 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_19) begin // @[Reg.scala 16:19]
      regData_r_4 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_23) begin // @[Reg.scala 16:19]
      regData_r_5 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_27) begin // @[Reg.scala 16:19]
      regData_r_6 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_31) begin // @[Reg.scala 16:19]
      regData_r_7 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_35) begin // @[Reg.scala 16:19]
      regData_r_8 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_39) begin // @[Reg.scala 16:19]
      regData_r_9 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_43) begin // @[Reg.scala 16:19]
      regData_r_10 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_47) begin // @[Reg.scala 16:19]
      regData_r_11 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_51) begin // @[Reg.scala 16:19]
      regData_r_12 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_55) begin // @[Reg.scala 16:19]
      regData_r_13 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_59) begin // @[Reg.scala 16:19]
      regData_r_14 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_63) begin // @[Reg.scala 16:19]
      regData_r_15 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_67) begin // @[Reg.scala 16:19]
      regData_r_16 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_71) begin // @[Reg.scala 16:19]
      regData_r_17 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_75) begin // @[Reg.scala 16:19]
      regData_r_18 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_79) begin // @[Reg.scala 16:19]
      regData_r_19 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_83) begin // @[Reg.scala 16:19]
      regData_r_20 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_87) begin // @[Reg.scala 16:19]
      regData_r_21 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_91) begin // @[Reg.scala 16:19]
      regData_r_22 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_95) begin // @[Reg.scala 16:19]
      regData_r_23 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_99) begin // @[Reg.scala 16:19]
      regData_r_24 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_103) begin // @[Reg.scala 16:19]
      regData_r_25 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_107) begin // @[Reg.scala 16:19]
      regData_r_26 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_111) begin // @[Reg.scala 16:19]
      regData_r_27 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_115) begin // @[Reg.scala 16:19]
      regData_r_28 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_119) begin // @[Reg.scala 16:19]
      regData_r_29 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_123) begin // @[Reg.scala 16:19]
      regData_r_30 <= io_din; // @[Reg.scala 16:23]
    end
    if (_regData_T_127) begin // @[Reg.scala 16:19]
      regData_r_31 <= io_din; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regData_r_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regData_r_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regData_r_3 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regData_r_4 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regData_r_5 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regData_r_6 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regData_r_7 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regData_r_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regData_r_9 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regData_r_10 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regData_r_11 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regData_r_12 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regData_r_13 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regData_r_14 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regData_r_15 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regData_r_16 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regData_r_17 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regData_r_18 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regData_r_19 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regData_r_20 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regData_r_21 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regData_r_22 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regData_r_23 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regData_r_24 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regData_r_25 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regData_r_26 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regData_r_27 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regData_r_28 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regData_r_29 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regData_r_30 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regData_r_31 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module iDecode(
  input         clock,
  input  [31:0] io_pc,
  input  [31:0] io_inst,
  input         io_regEn,
  output [63:0] io_dataEx_imme,
  output [63:0] io_dataEx_dOut1,
  output [63:0] io_dataEx_dOut2,
  input  [63:0] io_dataEx_dIn,
  output [63:0] io_dataEx_rdDout,
  output [4:0]  io_rdOut,
  input  [4:0]  io_rdIn,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  input  [4:0]  io_rsWB,
  output [63:0] io_dOutWB,
  input         block1,
  input         block23
);
  wire [31:0] imme_io_inst; // @[iDecode.scala 28:19]
  wire [63:0] imme_io_imme; // @[iDecode.scala 28:19]
  wire  rf_clock; // @[iDecode.scala 42:18]
  wire [31:0] rf_io_pc; // @[iDecode.scala 42:18]
  wire  rf_io_we; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs1; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rs2; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rd; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rdID; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout1; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_dout2; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_rdDout; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_din; // @[iDecode.scala 42:18]
  wire [4:0] rf_io_rsWB; // @[iDecode.scala 42:18]
  wire [63:0] rf_io_doutWB; // @[iDecode.scala 42:18]
  wire  rf_block1_0; // @[iDecode.scala 42:18]
  wire  rf_block23_0; // @[iDecode.scala 42:18]
  immeGen imme ( // @[iDecode.scala 28:19]
    .io_inst(imme_io_inst),
    .io_imme(imme_io_imme)
  );
  RF rf ( // @[iDecode.scala 42:18]
    .clock(rf_clock),
    .io_pc(rf_io_pc),
    .io_we(rf_io_we),
    .io_rs1(rf_io_rs1),
    .io_rs2(rf_io_rs2),
    .io_rd(rf_io_rd),
    .io_rdID(rf_io_rdID),
    .io_dout1(rf_io_dout1),
    .io_dout2(rf_io_dout2),
    .io_rdDout(rf_io_rdDout),
    .io_din(rf_io_din),
    .io_rsWB(rf_io_rsWB),
    .io_doutWB(rf_io_doutWB),
    .block1_0(rf_block1_0),
    .block23_0(rf_block23_0)
  );
  assign io_dataEx_imme = imme_io_imme; // @[iDecode.scala 30:18]
  assign io_dataEx_dOut1 = rf_io_dout1; // @[iDecode.scala 48:19]
  assign io_dataEx_dOut2 = rf_io_dout2; // @[iDecode.scala 49:19]
  assign io_dataEx_rdDout = rf_io_rdDout; // @[iDecode.scala 51:20]
  assign io_rdOut = io_inst[11:7]; // @[instDe.scala 20:16]
  assign io_rs1 = io_inst[19:15]; // @[instDe.scala 23:16]
  assign io_rs2 = io_inst[24:20]; // @[instDe.scala 26:16]
  assign io_dOutWB = rf_io_doutWB; // @[iDecode.scala 56:13]
  assign imme_io_inst = io_inst; // @[iDecode.scala 29:16]
  assign rf_clock = clock;
  assign rf_io_pc = io_pc; // @[iDecode.scala 53:12]
  assign rf_io_we = io_regEn; // @[iDecode.scala 46:12]
  assign rf_io_rs1 = io_inst[19:15]; // @[instDe.scala 23:16]
  assign rf_io_rs2 = io_inst[24:20]; // @[instDe.scala 26:16]
  assign rf_io_rd = io_rdIn; // @[iDecode.scala 45:12]
  assign rf_io_rdID = io_inst[11:7]; // @[instDe.scala 20:16]
  assign rf_io_din = io_dataEx_dIn; // @[iDecode.scala 47:13]
  assign rf_io_rsWB = io_rsWB; // @[iDecode.scala 55:14]
  assign rf_block1_0 = block1;
  assign rf_block23_0 = block23;
endmodule
module add(
  input         io_cin,
  input  [63:0] io_a,
  input  [63:0] io_b,
  output [63:0] io_sum,
  output        io_cout
);
  wire [64:0] _res_T = {1'h0,io_a}; // @[Cat.scala 30:58]
  wire [64:0] _res_T_1 = {1'h0,io_b}; // @[Cat.scala 30:58]
  wire [64:0] _res_T_3 = _res_T + _res_T_1; // @[add.scala 17:31]
  wire [64:0] _GEN_0 = {{64'd0}, io_cin}; // @[add.scala 17:52]
  wire [64:0] res = _res_T_3 + _GEN_0; // @[add.scala 17:52]
  assign io_sum = res[63:0]; // @[add.scala 18:18]
  assign io_cout = res[64]; // @[add.scala 19:19]
endmodule
module divR2(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_divw,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _dividend64Real_T_1 = io_dividend[63] & io_div_signed; // @[divR2.scala 21:51]
  wire [63:0] _dividend64Real_T_2 = ~io_dividend; // @[divR2.scala 21:70]
  wire [63:0] _dividend64Real_T_4 = _dividend64Real_T_2 + 64'h1; // @[divR2.scala 21:91]
  wire [63:0] dividend64Real = io_dividend[63] & io_div_signed ? _dividend64Real_T_4 : io_dividend; // @[divR2.scala 21:27]
  wire [63:0] _divisor64Real_T_2 = ~io_divisor; // @[divR2.scala 22:68]
  wire [63:0] _divisor64Real_T_4 = _divisor64Real_T_2 + 64'h1; // @[divR2.scala 22:88]
  wire [63:0] divisor64Real = io_divisor[63] & io_div_signed ? _divisor64Real_T_4 : io_divisor; // @[divR2.scala 22:26]
  wire  quoSgn64 = (io_dividend[63] ^ io_divisor[63]) & io_div_signed; // @[divR2.scala 23:67]
  wire  _dividend32Real_T_1 = io_dividend[31] & io_div_signed; // @[divR2.scala 26:48]
  wire [31:0] _dividend32Real_T_3 = ~io_dividend[31:0]; // @[divR2.scala 26:67]
  wire [31:0] _dividend32Real_T_5 = _dividend32Real_T_3 + 32'h1; // @[divR2.scala 26:94]
  wire [31:0] dividend32Real = io_dividend[31] & io_div_signed ? _dividend32Real_T_5 : io_dividend[31:0]; // @[divR2.scala 26:27]
  wire [31:0] _divisor32Real_T_3 = ~io_divisor[31:0]; // @[divR2.scala 27:65]
  wire [31:0] _divisor32Real_T_5 = _divisor32Real_T_3 + 32'h1; // @[divR2.scala 27:91]
  wire [31:0] divisor32Real = io_divisor[31] & io_div_signed ? _divisor32Real_T_5 : io_divisor[31:0]; // @[divR2.scala 27:26]
  wire  quoSgn32 = (io_dividend[31] ^ io_divisor[31]) & io_div_signed; // @[divR2.scala 28:61]
  reg [1:0] stateReg; // @[divR2.scala 35:25]
  wire  isDiv32 = stateReg == 2'h1; // @[divR2.scala 37:25]
  wire  isDiv64 = stateReg == 2'h2; // @[divR2.scala 38:26]
  reg [5:0] cnt; // @[divR2.scala 40:20]
  wire [1:0] _idleMux_T = {io_div_valid,io_divw}; // @[Cat.scala 30:58]
  wire [1:0] _idleMux_T_2 = 2'h3 == _idleMux_T ? 2'h1 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] idleMux = 2'h2 == _idleMux_T ? 2'h2 : _idleMux_T_2; // @[Mux.scala 80:57]
  wire [1:0] div32Mux = cnt == 6'h1f ? 2'h3 : 2'h1; // @[divR2.scala 49:21]
  wire [5:0] _cnt_T_2 = cnt + 6'h1; // @[divR2.scala 63:38]
  reg [127:0] dividendReg; // @[divR2.scala 66:28]
  reg [63:0] resReg; // @[divR2.scala 67:23]
  wire [127:0] _idleDividendMux_T_1 = {96'h0,dividend32Real}; // @[Cat.scala 30:58]
  wire [127:0] _idleDividendMux_T_2 = {64'h0,dividend64Real}; // @[Cat.scala 30:58]
  wire [127:0] _idleDividendMux_T_4 = 2'h3 == _idleMux_T ? _idleDividendMux_T_1 : 128'h0; // @[Mux.scala 80:57]
  wire [127:0] idleDividendMux = 2'h2 == _idleMux_T ? _idleDividendMux_T_2 : _idleDividendMux_T_4; // @[Mux.scala 80:57]
  wire [30:0] div32DividendMux_lo_hi = dividendReg[30:0]; // @[divR2.scala 78:59]
  wire [32:0] subed32 = dividendReg[63:31]; // @[divR2.scala 95:27]
  wire [32:0] _GEN_0 = {{1'd0}, divisor32Real}; // @[divR2.scala 96:26]
  wire [32:0] subRes32 = subed32 - _GEN_0; // @[divR2.scala 96:26]
  wire [31:0] rem32M = subRes32[32] ? subed32[31:0] : subRes32[31:0]; // @[divR2.scala 97:16]
  wire [127:0] div32DividendMux = {64'h0,rem32M,div32DividendMux_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [62:0] div64DividendMux_hi_lo = dividendReg[62:0]; // @[divR2.scala 79:48]
  wire [64:0] subed64 = dividendReg[127:63]; // @[divR2.scala 91:29]
  wire [64:0] _GEN_1 = {{1'd0}, divisor64Real}; // @[divR2.scala 92:26]
  wire [64:0] subRes64 = subed64 - _GEN_1; // @[divR2.scala 92:26]
  wire [63:0] rem64M = subRes64[64] ? subed64[63:0] : subRes64[63:0]; // @[divR2.scala 93:16]
  wire [127:0] div64DividendMux = {rem64M,div64DividendMux_hi_lo,1'h0}; // @[Cat.scala 30:58]
  wire [62:0] resReg_hi = resReg[62:0]; // @[divR2.scala 104:31]
  wire  resReg_lo = ~subRes32[32]; // @[divR2.scala 104:38]
  wire [63:0] _resReg_T_1 = {resReg_hi,resReg_lo}; // @[Cat.scala 30:58]
  wire  resReg_lo_1 = ~subRes64[64]; // @[divR2.scala 105:38]
  wire [63:0] _resReg_T_3 = {resReg_hi,resReg_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _res64Out_T = ~resReg; // @[divR2.scala 110:35]
  wire [63:0] _res64Out_T_2 = _res64Out_T + 64'h1; // @[divR2.scala 110:53]
  wire [63:0] res64Out = quoSgn64 ? _res64Out_T_2 : resReg; // @[divR2.scala 110:21]
  wire [63:0] _rem64Out_T_1 = ~dividendReg[127:64]; // @[divR2.scala 111:32]
  wire [63:0] _rem64Out_T_3 = _rem64Out_T_1 + 64'h1; // @[divR2.scala 111:63]
  wire [63:0] rem64Out = _dividend64Real_T_1 ? _rem64Out_T_3 : dividendReg[127:64]; // @[divR2.scala 111:20]
  wire [31:0] _res32out_T_1 = ~resReg[31:0]; // @[divR2.scala 113:56]
  wire [31:0] res32out_lo = _res32out_T_1 + 32'h1; // @[divR2.scala 113:79]
  wire [63:0] _res32out_T_3 = {32'hffffffff,res32out_lo}; // @[Cat.scala 30:58]
  wire [63:0] res32out = quoSgn32 ? _res32out_T_3 : resReg; // @[divR2.scala 113:21]
  wire [31:0] _rem32Out_T_1 = ~dividendReg[63:32]; // @[divR2.scala 115:56]
  wire [31:0] rem32Out_lo = _rem32Out_T_1 + 32'h1; // @[divR2.scala 115:85]
  wire [63:0] _rem32Out_T_3 = {32'hffffffff,rem32Out_lo}; // @[Cat.scala 30:58]
  wire [63:0] _rem32Out_T_4 = {32'h0,dividendReg[63:32]}; // @[Cat.scala 30:58]
  wire [63:0] rem32Out = _dividend32Real_T_1 ? _rem32Out_T_3 : _rem32Out_T_4; // @[divR2.scala 115:21]
  assign io_out_valid = stateReg == 2'h3; // @[divR2.scala 39:27]
  assign io_quotient = io_divw ? res32out : res64Out; // @[divR2.scala 119:21]
  assign io_remainder = io_divw ? rem32Out : rem64Out; // @[divR2.scala 120:22]
  always @(posedge clock) begin
    if (reset) begin // @[divR2.scala 35:25]
      stateReg <= 2'h0; // @[divR2.scala 35:25]
    end else if (2'h3 == stateReg) begin // @[Mux.scala 80:57]
      if (io_block) begin // @[divR2.scala 51:22]
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h0;
      end
    end else if (2'h2 == stateReg) begin // @[Mux.scala 80:57]
      if (cnt == 6'h3f) begin // @[divR2.scala 50:21]
        stateReg <= 2'h3;
      end else begin
        stateReg <= 2'h2;
      end
    end else if (2'h1 == stateReg) begin // @[Mux.scala 80:57]
      stateReg <= div32Mux;
    end else begin
      stateReg <= idleMux;
    end
    if (reset) begin // @[divR2.scala 40:20]
      cnt <= 6'h0; // @[divR2.scala 40:20]
    end else if (isDiv32 | isDiv64) begin // @[divR2.scala 63:13]
      cnt <= _cnt_T_2;
    end else begin
      cnt <= 6'h0;
    end
    if (reset) begin // @[divR2.scala 66:28]
      dividendReg <= 128'h0; // @[divR2.scala 66:28]
    end else if (!(2'h3 == stateReg)) begin // @[Mux.scala 80:57]
      if (2'h2 == stateReg) begin // @[Mux.scala 80:57]
        dividendReg <= div64DividendMux;
      end else if (2'h1 == stateReg) begin // @[Mux.scala 80:57]
        dividendReg <= div32DividendMux;
      end else begin
        dividendReg <= idleDividendMux;
      end
    end
    if (reset) begin // @[divR2.scala 67:23]
      resReg <= 64'h0; // @[divR2.scala 67:23]
    end else if (!(2'h3 == stateReg)) begin // @[Mux.scala 80:57]
      if (2'h2 == stateReg) begin // @[Mux.scala 80:57]
        resReg <= _resReg_T_3;
      end else if (2'h1 == stateReg) begin // @[Mux.scala 80:57]
        resReg <= _resReg_T_1;
      end else begin
        resReg <= 64'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {4{`RANDOM}};
  dividendReg = _RAND_2[127:0];
  _RAND_3 = {2{`RANDOM}};
  resReg = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module boothSel(
  input  [2:0]   io_y,
  input  [131:0] io_x,
  output [131:0] io_p,
  output         io_c
);
  wire  _selNegative_T_3 = ~io_y[0]; // @[mul.scala 13:42]
  wire  _selNegative_T_6 = ~io_y[1]; // @[mul.scala 13:53]
  wire  _selNegative_T_9 = io_y[1] & ~io_y[0] | ~io_y[1] & io_y[0]; // @[mul.scala 13:51]
  wire  selNegative = io_y[2] & (io_y[1] & ~io_y[0] | ~io_y[1] & io_y[0]); // @[mul.scala 13:29]
  wire  _selPositive_T_1 = ~io_y[2]; // @[mul.scala 14:21]
  wire  selPositive = ~io_y[2] & _selNegative_T_9; // @[mul.scala 14:30]
  wire  selDoubleNegative = io_y[2] & _selNegative_T_6 & _selNegative_T_3; // @[mul.scala 15:46]
  wire  selDoublePositive = _selPositive_T_1 & io_y[1] & io_y[0]; // @[mul.scala 16:46]
  wire [131:0] _io_p_T_1 = selNegative ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _io_p_T_2 = ~io_x; // @[mul.scala 18:42]
  wire [131:0] _io_p_T_3 = _io_p_T_1 & _io_p_T_2; // @[mul.scala 18:39]
  wire [131:0] _io_p_T_5 = selDoubleNegative ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [130:0] io_p_hi = ~io_x[130:0]; // @[mul.scala 19:50]
  wire [131:0] _io_p_T_7 = {io_p_hi,1'h1}; // @[Cat.scala 30:58]
  wire [131:0] _io_p_T_8 = _io_p_T_5 & _io_p_T_7; // @[mul.scala 19:45]
  wire [131:0] _io_p_T_9 = _io_p_T_3 | _io_p_T_8; // @[mul.scala 18:56]
  wire [131:0] _io_p_T_11 = selPositive ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _io_p_T_12 = _io_p_T_11 & io_x; // @[mul.scala 20:39]
  wire [131:0] _io_p_T_13 = _io_p_T_9 | _io_p_T_12; // @[mul.scala 19:79]
  wire [131:0] _io_p_T_15 = selDoublePositive ? 132'hfffffffffffffffffffffffffffffffff : 132'h0; // @[Bitwise.scala 72:12]
  wire [131:0] _io_p_T_16 = {io_x[130:0],1'h0}; // @[Cat.scala 30:58]
  wire [131:0] _io_p_T_17 = _io_p_T_15 & _io_p_T_16; // @[mul.scala 21:46]
  assign io_p = _io_p_T_13 | _io_p_T_17; // @[mul.scala 20:45]
  assign io_c = selDoubleNegative | selNegative; // @[mul.scala 23:29]
endmodule
module add_1(
  input          io_cin,
  input  [131:0] io_a,
  input  [131:0] io_b,
  output [131:0] io_sum
);
  wire [132:0] _res_T = {1'h0,io_a}; // @[Cat.scala 30:58]
  wire [132:0] _res_T_1 = {1'h0,io_b}; // @[Cat.scala 30:58]
  wire [132:0] _res_T_3 = _res_T + _res_T_1; // @[add.scala 17:31]
  wire [132:0] _GEN_0 = {{132'd0}, io_cin}; // @[add.scala 17:52]
  wire [132:0] res = _res_T_3 + _GEN_0; // @[add.scala 17:52]
  assign io_sum = res[131:0]; // @[add.scala 18:18]
endmodule
module mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [63:0] io_result_low,
  input         io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] boothIns_io_y; // @[mul.scala 103:24]
  wire [131:0] boothIns_io_x; // @[mul.scala 103:24]
  wire [131:0] boothIns_io_p; // @[mul.scala 103:24]
  wire  boothIns_io_c; // @[mul.scala 103:24]
  wire  addIns_io_cin; // @[mul.scala 105:22]
  wire [131:0] addIns_io_a; // @[mul.scala 105:22]
  wire [131:0] addIns_io_b; // @[mul.scala 105:22]
  wire [131:0] addIns_io_sum; // @[mul.scala 105:22]
  reg [1:0] stateReg; // @[mul.scala 40:25]
  wire  isIdle = stateReg == 2'h0; // @[mul.scala 41:25]
  wire  isMul = stateReg == 2'h1; // @[mul.scala 42:24]
  reg [5:0] cnt; // @[mul.scala 47:20]
  wire [1:0] idleMux = io_mul_valid ? 2'h1 : 2'h0; // @[mul.scala 53:20]
  wire [5:0] _cnt_T_1 = cnt + 6'h1; // @[mul.scala 65:25]
  wire [66:0] multiplierEx = {2'h0,io_multiplier,1'h0}; // @[Cat.scala 30:58]
  reg [66:0] multiplierReg; // @[mul.scala 80:30]
  wire  _multiplierReg_T = isIdle & io_mul_valid; // @[mul.scala 82:12]
  wire [64:0] multiplierReg_lo = multiplierReg[66:2]; // @[mul.scala 86:34]
  wire [66:0] _multiplierReg_T_1 = {2'h0,multiplierReg_lo}; // @[Cat.scala 30:58]
  reg [131:0] multiplicandReg; // @[mul.scala 91:32]
  wire [131:0] _multiplicandReg_T_1 = {66'h0,2'h0,io_multiplicand}; // @[Cat.scala 30:58]
  wire [129:0] multiplicandReg_hi = multiplicandReg[129:0]; // @[mul.scala 97:26]
  wire [131:0] _multiplicandReg_T_2 = {multiplicandReg_hi,2'h0}; // @[Cat.scala 30:58]
  reg [131:0] resReg; // @[mul.scala 104:23]
  boothSel boothIns ( // @[mul.scala 103:24]
    .io_y(boothIns_io_y),
    .io_x(boothIns_io_x),
    .io_p(boothIns_io_p),
    .io_c(boothIns_io_c)
  );
  add_1 addIns ( // @[mul.scala 105:22]
    .io_cin(addIns_io_cin),
    .io_a(addIns_io_a),
    .io_b(addIns_io_b),
    .io_sum(addIns_io_sum)
  );
  assign io_out_valid = stateReg == 2'h2; // @[mul.scala 43:24]
  assign io_result_low = resReg[63:0]; // @[mul.scala 137:26]
  assign boothIns_io_y = multiplierReg[2:0]; // @[mul.scala 107:32]
  assign boothIns_io_x = multiplicandReg; // @[mul.scala 108:16]
  assign addIns_io_cin = boothIns_io_c; // @[mul.scala 111:17]
  assign addIns_io_a = boothIns_io_p; // @[mul.scala 110:15]
  assign addIns_io_b = resReg; // @[mul.scala 112:15]
  always @(posedge clock) begin
    if (reset) begin // @[mul.scala 40:25]
      stateReg <= 2'h0; // @[mul.scala 40:25]
    end else if (2'h2 == stateReg) begin // @[Mux.scala 80:57]
      if (io_block) begin // @[mul.scala 55:22]
        stateReg <= 2'h2;
      end else begin
        stateReg <= 2'h0;
      end
    end else if (2'h1 == stateReg) begin // @[Mux.scala 80:57]
      if (cnt == 6'h20) begin // @[mul.scala 54:19]
        stateReg <= 2'h2;
      end else begin
        stateReg <= 2'h1;
      end
    end else if (2'h0 == stateReg) begin // @[Mux.scala 80:57]
      stateReg <= idleMux;
    end else begin
      stateReg <= 2'h0;
    end
    if (reset) begin // @[mul.scala 47:20]
      cnt <= 6'h0; // @[mul.scala 47:20]
    end else if (isMul) begin // @[mul.scala 65:13]
      cnt <= _cnt_T_1;
    end else begin
      cnt <= 6'h0;
    end
    if (reset) begin // @[mul.scala 80:30]
      multiplierReg <= 67'h0; // @[mul.scala 80:30]
    end else if (_multiplierReg_T) begin // @[mul.scala 81:23]
      multiplierReg <= multiplierEx;
    end else if (isMul) begin // @[mul.scala 84:8]
      multiplierReg <= _multiplierReg_T_1;
    end
    if (reset) begin // @[mul.scala 91:32]
      multiplicandReg <= 132'h0; // @[mul.scala 91:32]
    end else if (_multiplierReg_T) begin // @[mul.scala 92:25]
      multiplicandReg <= _multiplicandReg_T_1;
    end else if (isMul) begin // @[mul.scala 95:8]
      multiplicandReg <= _multiplicandReg_T_2;
    end
    if (reset) begin // @[mul.scala 104:23]
      resReg <= 132'h0; // @[mul.scala 104:23]
    end else if (isIdle) begin // @[mul.scala 117:16]
      resReg <= 132'h0;
    end else if (isMul) begin // @[mul.scala 120:8]
      resReg <= addIns_io_sum;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {3{`RANDOM}};
  multiplierReg = _RAND_2[66:0];
  _RAND_3 = {5{`RANDOM}};
  multiplicandReg = _RAND_3[131:0];
  _RAND_4 = {5{`RANDOM}};
  resReg = _RAND_4[131:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_srcA,
  input  [63:0] io_srcB,
  input  [4:0]  io_ALUCtrl,
  output [63:0] io_ALUResult,
  output        block1_0,
  input         block23_0
);
  wire  addIns_io_cin; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_a; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_b; // @[ALU.scala 21:22]
  wire [63:0] addIns_io_sum; // @[ALU.scala 21:22]
  wire  addIns_io_cout; // @[ALU.scala 21:22]
  wire  divR2Ins_clock; // @[ALU.scala 31:23]
  wire  divR2Ins_reset; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_dividend; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_divisor; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_valid; // @[ALU.scala 31:23]
  wire  divR2Ins_io_divw; // @[ALU.scala 31:23]
  wire  divR2Ins_io_div_signed; // @[ALU.scala 31:23]
  wire  divR2Ins_io_out_valid; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_quotient; // @[ALU.scala 31:23]
  wire [63:0] divR2Ins_io_remainder; // @[ALU.scala 31:23]
  wire  divR2Ins_io_block; // @[ALU.scala 31:23]
  wire  mulIns_clock; // @[ALU.scala 46:22]
  wire  mulIns_reset; // @[ALU.scala 46:22]
  wire  mulIns_io_mul_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplicand; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_multiplier; // @[ALU.scala 46:22]
  wire  mulIns_io_out_valid; // @[ALU.scala 46:22]
  wire [63:0] mulIns_io_result_low; // @[ALU.scala 46:22]
  wire  mulIns_io_block; // @[ALU.scala 46:22]
  wire  sub = io_ALUCtrl == 5'h1 | io_ALUCtrl == 5'h5 | io_ALUCtrl == 5'h10 | io_ALUCtrl == 5'h5 | io_ALUCtrl == 5'h7 |
    io_ALUCtrl == 5'h1b | io_ALUCtrl == 5'h1c; // @[ALU.scala 23:56]
  wire [63:0] srcBInv = ~io_srcB; // @[ALU.scala 24:18]
  wire  _divValid_T_4 = io_ALUCtrl == 5'h14; // @[ALU.scala 33:79]
  wire  _divValid_T_5 = io_ALUCtrl == 5'h11 | io_ALUCtrl == 5'h12 | io_ALUCtrl == 5'h14; // @[ALU.scala 33:66]
  wire  _divValid_T_6 = io_ALUCtrl == 5'h15; // @[ALU.scala 33:79]
  wire  _divValid_T_10 = io_ALUCtrl == 5'h18; // @[ALU.scala 33:79]
  wire  _divValid_T_12 = io_ALUCtrl == 5'h19; // @[ALU.scala 33:79]
  wire [31:0] srcAUSignW_lo = io_srcA[31:0]; // @[ALU.scala 47:35]
  wire [63:0] srcAUSignW = {32'h0,srcAUSignW_lo}; // @[Cat.scala 30:58]
  wire [31:0] srcBUSignW_lo = io_srcB[31:0]; // @[ALU.scala 48:35]
  wire [63:0] srcBUSignW = {32'h0,srcBUSignW_lo}; // @[Cat.scala 30:58]
  wire  _mulValid_T = io_ALUCtrl == 5'h13; // @[ALU.scala 50:79]
  wire [5:0] shamt = io_srcB[5:0]; // @[ALU.scala 61:22]
  wire [63:0] _T_2 = $signed(io_srcA) >>> shamt; // @[ALU.scala 65:42]
  wire [63:0] _T_3 = io_srcA >> shamt; // @[ALU.scala 66:25]
  wire [126:0] _GEN_0 = {{63'd0}, io_srcA}; // @[ALU.scala 67:25]
  wire [126:0] _T_4 = _GEN_0 << shamt; // @[ALU.scala 67:25]
  wire  _T_6 = ~addIns_io_cout; // @[ALU.scala 69:16]
  wire [63:0] _T_7 = io_srcA & io_srcB; // @[ALU.scala 70:25]
  wire [63:0] _T_8 = io_srcA | io_srcB; // @[ALU.scala 71:24]
  wire [63:0] _T_9 = io_srcA ^ io_srcB; // @[ALU.scala 72:25]
  wire  lo = io_srcA != io_srcB; // @[ALU.scala 73:32]
  wire [63:0] _T_10 = {63'h0,lo}; // @[Cat.scala 30:58]
  wire [31:0] lo_1 = srcAUSignW_lo >> shamt; // @[ALU.scala 74:48]
  wire  signBit = lo_1[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi = signBit ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_13 = {hi,lo_1}; // @[Cat.scala 30:58]
  wire [31:0] lo_2 = addIns_io_sum[31:0]; // @[ALU.scala 75:40]
  wire  signBit_1 = lo_2[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_1 = signBit_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {hi_1,lo_2}; // @[Cat.scala 30:58]
  wire [94:0] _GEN_1 = {{63'd0}, srcAUSignW_lo}; // @[ALU.scala 76:48]
  wire [94:0] _T_17 = _GEN_1 << shamt; // @[ALU.scala 76:48]
  wire [31:0] lo_3 = _T_17[31:0]; // @[ALU.scala 76:58]
  wire  signBit_2 = lo_3[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_2 = signBit_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_19 = {hi_2,lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _T_21 = io_srcA[31:0]; // @[ALU.scala 77:41]
  wire [31:0] lo_4 = $signed(_T_21) >>> shamt; // @[ALU.scala 77:65]
  wire  signBit_3 = lo_4[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_3 = signBit_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_24 = {hi_3,lo_4}; // @[Cat.scala 30:58]
  wire [31:0] lo_6 = divR2Ins_io_quotient[31:0]; // @[ALU.scala 79:46]
  wire  signBit_5 = lo_6[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_5 = signBit_5 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_28 = {hi_5,lo_6}; // @[Cat.scala 30:58]
  wire [31:0] lo_7 = divR2Ins_io_remainder[31:0]; // @[ALU.scala 80:47]
  wire  signBit_6 = lo_7[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_6 = signBit_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_30 = {hi_6,lo_7}; // @[Cat.scala 30:58]
  wire [31:0] lo_8 = mulIns_io_result_low[31:0]; // @[ALU.scala 81:45]
  wire  signBit_7 = lo_8[31]; // @[immeGen.scala 17:22]
  wire [31:0] hi_7 = signBit_7 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_32 = {hi_7,lo_8}; // @[Cat.scala 30:58]
  wire  _T_37 = io_srcA == io_srcB; // @[ALU.scala 88:24]
  wire  _T_39 = ~addIns_io_sum[63]; // @[ALU.scala 91:16]
  wire [63:0] _io_ALUResult_T_1 = 5'h0 == io_ALUCtrl ? addIns_io_sum : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_ALUResult_T_3 = 5'h1 == io_ALUCtrl ? addIns_io_sum : _io_ALUResult_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_ALUResult_T_5 = 5'h9 == io_ALUCtrl ? _T_2 : _io_ALUResult_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_ALUResult_T_7 = 5'h8 == io_ALUCtrl ? _T_3 : _io_ALUResult_T_5; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_9 = 5'h6 == io_ALUCtrl ? _T_4 : {{63'd0}, _io_ALUResult_T_7}; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_11 = 5'h5 == io_ALUCtrl ? {{126'd0}, addIns_io_sum[63]} : _io_ALUResult_T_9; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_13 = 5'h7 == io_ALUCtrl ? {{126'd0}, _T_6} : _io_ALUResult_T_11; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_15 = 5'h2 == io_ALUCtrl ? {{63'd0}, _T_7} : _io_ALUResult_T_13; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_17 = 5'h3 == io_ALUCtrl ? {{63'd0}, _T_8} : _io_ALUResult_T_15; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_19 = 5'h4 == io_ALUCtrl ? {{63'd0}, _T_9} : _io_ALUResult_T_17; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_21 = 5'hb == io_ALUCtrl ? {{63'd0}, _T_10} : _io_ALUResult_T_19; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_23 = 5'hc == io_ALUCtrl ? {{63'd0}, _T_13} : _io_ALUResult_T_21; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_25 = 5'hd == io_ALUCtrl ? {{63'd0}, _T_15} : _io_ALUResult_T_23; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_27 = 5'he == io_ALUCtrl ? {{63'd0}, _T_19} : _io_ALUResult_T_25; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_29 = 5'hf == io_ALUCtrl ? {{63'd0}, _T_24} : _io_ALUResult_T_27; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_31 = 5'h10 == io_ALUCtrl ? {{63'd0}, _T_15} : _io_ALUResult_T_29; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_33 = 5'h11 == io_ALUCtrl ? {{63'd0}, _T_28} : _io_ALUResult_T_31; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_35 = 5'h12 == io_ALUCtrl ? {{63'd0}, _T_30} : _io_ALUResult_T_33; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_37 = 5'h13 == io_ALUCtrl ? {{63'd0}, _T_32} : _io_ALUResult_T_35; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_39 = 5'h14 == io_ALUCtrl ? {{63'd0}, _T_30} : _io_ALUResult_T_37; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_41 = 5'h15 == io_ALUCtrl ? {{63'd0}, _T_28} : _io_ALUResult_T_39; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_43 = 5'h16 == io_ALUCtrl ? {{63'd0}, mulIns_io_result_low} : _io_ALUResult_T_41; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_45 = 5'h17 == io_ALUCtrl ? {{63'd0}, divR2Ins_io_quotient} : _io_ALUResult_T_43; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_47 = 5'h18 == io_ALUCtrl ? {{63'd0}, divR2Ins_io_remainder} : _io_ALUResult_T_45; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_49 = 5'h19 == io_ALUCtrl ? {{63'd0}, divR2Ins_io_quotient} : _io_ALUResult_T_47; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_51 = 5'h1a == io_ALUCtrl ? {{126'd0}, _T_37} : _io_ALUResult_T_49; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_53 = 5'h1b == io_ALUCtrl ? {{126'd0}, addIns_io_cout} : _io_ALUResult_T_51; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_55 = 5'h1c == io_ALUCtrl ? {{126'd0}, _T_39} : _io_ALUResult_T_53; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_57 = 5'h1d == io_ALUCtrl ? {{63'd0}, divR2Ins_io_remainder} : _io_ALUResult_T_55; // @[Mux.scala 80:57]
  wire [126:0] _io_ALUResult_T_59 = 5'ha == io_ALUCtrl ? {{63'd0}, io_srcA} : _io_ALUResult_T_57; // @[Mux.scala 80:57]
  wire  block1 = divR2Ins_io_div_valid & ~divR2Ins_io_out_valid | mulIns_io_mul_valid & ~mulIns_io_out_valid; // @[ALU.scala 98:61]
  add addIns ( // @[ALU.scala 21:22]
    .io_cin(addIns_io_cin),
    .io_a(addIns_io_a),
    .io_b(addIns_io_b),
    .io_sum(addIns_io_sum),
    .io_cout(addIns_io_cout)
  );
  divR2 divR2Ins ( // @[ALU.scala 31:23]
    .clock(divR2Ins_clock),
    .reset(divR2Ins_reset),
    .io_dividend(divR2Ins_io_dividend),
    .io_divisor(divR2Ins_io_divisor),
    .io_div_valid(divR2Ins_io_div_valid),
    .io_divw(divR2Ins_io_divw),
    .io_div_signed(divR2Ins_io_div_signed),
    .io_out_valid(divR2Ins_io_out_valid),
    .io_quotient(divR2Ins_io_quotient),
    .io_remainder(divR2Ins_io_remainder),
    .io_block(divR2Ins_io_block)
  );
  mul mulIns ( // @[ALU.scala 46:22]
    .clock(mulIns_clock),
    .reset(mulIns_reset),
    .io_mul_valid(mulIns_io_mul_valid),
    .io_multiplicand(mulIns_io_multiplicand),
    .io_multiplier(mulIns_io_multiplier),
    .io_out_valid(mulIns_io_out_valid),
    .io_result_low(mulIns_io_result_low),
    .io_block(mulIns_io_block)
  );
  assign io_ALUResult = _io_ALUResult_T_59[63:0]; // @[ALU.scala 95:16]
  assign block1_0 = block1;
  assign addIns_io_cin = io_ALUCtrl == 5'h1 | io_ALUCtrl == 5'h5 | io_ALUCtrl == 5'h10 | io_ALUCtrl == 5'h5 | io_ALUCtrl
     == 5'h7 | io_ALUCtrl == 5'h1b | io_ALUCtrl == 5'h1c; // @[ALU.scala 23:56]
  assign addIns_io_a = io_srcA; // @[ALU.scala 26:15]
  assign addIns_io_b = sub ? srcBInv : io_srcB; // @[ALU.scala 28:21]
  assign divR2Ins_clock = clock;
  assign divR2Ins_reset = reset;
  assign divR2Ins_io_dividend = io_srcA; // @[ALU.scala 38:24]
  assign divR2Ins_io_divisor = io_srcB; // @[ALU.scala 39:23]
  assign divR2Ins_io_div_valid = io_ALUCtrl == 5'h11 | io_ALUCtrl == 5'h12 | io_ALUCtrl == 5'h14 | io_ALUCtrl == 5'h15
     | io_ALUCtrl == 5'h17 | io_ALUCtrl == 5'h18 | io_ALUCtrl == 5'h19 | io_ALUCtrl == 5'h1d; // @[ALU.scala 33:66]
  assign divR2Ins_io_divw = _divValid_T_5 | _divValid_T_6; // @[ALU.scala 35:58]
  assign divR2Ins_io_div_signed = _divValid_T_4 | _divValid_T_6 | _divValid_T_10 | _divValid_T_12; // @[ALU.scala 37:68]
  assign divR2Ins_io_block = block23_0; // @[ALU.scala 105:21]
  assign mulIns_clock = clock;
  assign mulIns_reset = reset;
  assign mulIns_io_mul_valid = io_ALUCtrl == 5'h13 | io_ALUCtrl == 5'h16; // @[ALU.scala 50:66]
  assign mulIns_io_multiplicand = _mulValid_T ? srcAUSignW : io_srcA; // @[ALU.scala 56:32]
  assign mulIns_io_multiplier = _mulValid_T ? srcBUSignW : io_srcB; // @[ALU.scala 57:30]
  assign mulIns_io_block = block23_0; // @[ALU.scala 105:21]
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_csrrwen,
  input         io_csrswen,
  input         io_csrrsien,
  input         io_csrrcien,
  input         io_csrrcen,
  input         io_csrrwien,
  input         io_ecall,
  input  [63:0] io_rs1,
  input  [11:0] io_imme,
  input  [63:0] io_pc,
  input  [4:0]  io_uimm,
  output [63:0] io_rd,
  output [63:0] io_mtvec,
  output [63:0] io_mepc,
  input         io_mret,
  input         intrTimeCnt_0,
  output        startTimeCnt_0,
  input         blockDMA_0,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  intr = intrTimeCnt_0 & io_pc != 64'h0; // @[CSR.scala 37:26]
  wire  csren = io_csrrwen | io_csrswen | io_csrrcen | io_csrrsien | io_csrrcien | io_csrrwien; // @[CSR.scala 54:82]
  wire [5:0] sel1H = {io_csrrwien,io_csrrcien,io_csrrsien,io_csrrcen,io_csrswen,io_csrrwen}; // @[Cat.scala 30:58]
  wire [63:0] uimmext = {59'h0,io_uimm}; // @[Cat.scala 30:58]
  wire  mepcen = io_ecall | csren & io_imme == 12'h341 | intr; // @[CSR.scala 58:58]
  wire  _mepcval_T = io_ecall | intr; // @[CSR.scala 61:14]
  reg [63:0] mepcins_r; // @[Reg.scala 27:20]
  wire [63:0] _mepcval_T_1 = io_rs1 | mepcins_r; // @[CSR.scala 67:15]
  wire [63:0] _mepcval_T_2 = ~io_rs1; // @[CSR.scala 68:10]
  wire [63:0] _mepcval_T_3 = _mepcval_T_2 & mepcins_r; // @[CSR.scala 68:28]
  wire [63:0] _mepcval_T_4 = uimmext | mepcins_r; // @[CSR.scala 69:17]
  wire [63:0] _mepcval_T_5 = ~uimmext; // @[CSR.scala 70:10]
  wire [63:0] _mepcval_T_6 = _mepcval_T_5 & mepcins_r; // @[CSR.scala 70:29]
  wire [63:0] _mepcval_T_13 = sel1H[0] ? io_rs1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_14 = sel1H[1] ? _mepcval_T_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_15 = sel1H[2] ? _mepcval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_16 = sel1H[3] ? _mepcval_T_4 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_17 = sel1H[4] ? _mepcval_T_6 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_18 = sel1H[5] ? uimmext : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_19 = _mepcval_T_13 | _mepcval_T_14; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_20 = _mepcval_T_19 | _mepcval_T_15; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_21 = _mepcval_T_20 | _mepcval_T_16; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_22 = _mepcval_T_21 | _mepcval_T_17; // @[Mux.scala 27:72]
  wire [63:0] _mepcval_T_23 = _mepcval_T_22 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mepcins_T = block1_0 | block23_0; // @[CSR.scala 75:56]
  wire  _mepcins_T_2 = ~(block1_0 | block23_0 | blockDMA_0); // @[CSR.scala 75:47]
  wire  _mepcins_T_3 = mepcen & ~(block1_0 | block23_0 | blockDMA_0); // @[CSR.scala 75:44]
  wire  mcauseen = io_ecall | csren & io_imme == 12'h342 | intr; // @[CSR.scala 77:61]
  reg [63:0] mcauseins_r; // @[Reg.scala 27:20]
  wire [63:0] _mcauseval_T = io_rs1 | mcauseins_r; // @[CSR.scala 89:16]
  wire [63:0] _mcauseval_T_2 = _mepcval_T_2 & mcauseins_r; // @[CSR.scala 90:28]
  wire [63:0] _mcauseval_T_3 = uimmext | mcauseins_r; // @[CSR.scala 91:17]
  wire [63:0] _mcauseval_T_5 = _mepcval_T_5 & mcauseins_r; // @[CSR.scala 92:29]
  wire [63:0] _mcauseval_T_13 = sel1H[1] ? _mcauseval_T : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_14 = sel1H[2] ? _mcauseval_T_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_15 = sel1H[3] ? _mcauseval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_16 = sel1H[4] ? _mcauseval_T_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_18 = _mepcval_T_13 | _mcauseval_T_13; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_19 = _mcauseval_T_18 | _mcauseval_T_14; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_20 = _mcauseval_T_19 | _mcauseval_T_15; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_21 = _mcauseval_T_20 | _mcauseval_T_16; // @[Mux.scala 27:72]
  wire [63:0] _mcauseval_T_22 = _mcauseval_T_21 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mcauseins_T_3 = mcauseen & _mepcins_T_2; // @[CSR.scala 97:50]
  wire  mtvecen = csren & io_imme == 12'h305; // @[CSR.scala 99:25]
  reg [63:0] mtvecins_r; // @[Reg.scala 27:20]
  wire [63:0] _mtvecval_T = io_rs1 | mtvecins_r; // @[CSR.scala 105:14]
  wire [63:0] _mtvecval_T_2 = _mepcval_T_2 & mtvecins_r; // @[CSR.scala 106:26]
  wire [63:0] _mtvecval_T_3 = uimmext | mtvecins_r; // @[CSR.scala 107:15]
  wire [63:0] _mtvecval_T_5 = _mepcval_T_5 & mtvecins_r; // @[CSR.scala 108:27]
  wire [63:0] _mtvecval_T_13 = sel1H[1] ? _mtvecval_T : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_14 = sel1H[2] ? _mtvecval_T_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_15 = sel1H[3] ? _mtvecval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_16 = sel1H[4] ? _mtvecval_T_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_18 = _mepcval_T_13 | _mtvecval_T_13; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_19 = _mtvecval_T_18 | _mtvecval_T_14; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_20 = _mtvecval_T_19 | _mtvecval_T_15; // @[Mux.scala 27:72]
  wire [63:0] _mtvecval_T_21 = _mtvecval_T_20 | _mtvecval_T_16; // @[Mux.scala 27:72]
  wire [63:0] mtvecval = _mtvecval_T_21 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mtvecins_T_3 = ~(_mepcins_T | intr | blockDMA_0); // @[CSR.scala 112:50]
  wire  _mtvecins_T_4 = mtvecen & ~(_mepcins_T | intr | blockDMA_0); // @[CSR.scala 112:47]
  wire  mstatusen = csren & io_imme == 12'h300 | io_ecall | intr | io_mret; // @[CSR.scala 114:73]
  reg [63:0] mstatusins_r; // @[Reg.scala 27:20]
  wire [55:0] mstatusval_hi_hi_hi = mstatusins_r[63:8]; // @[CSR.scala 119:19]
  wire  mstatusval_hi_hi_lo = mstatusins_r[3]; // @[CSR.scala 119:44]
  wire [2:0] mstatusval_hi_lo = mstatusins_r[6:4]; // @[CSR.scala 119:58]
  wire [2:0] mstatusval_lo_lo = mstatusins_r[2:0]; // @[CSR.scala 119:82]
  wire [63:0] _mstatusval_T_1 = {mstatusval_hi_hi_hi,mstatusval_hi_hi_lo,mstatusval_hi_lo,1'h0,mstatusval_lo_lo}; // @[Cat.scala 30:58]
  wire  mstatusval_lo_hi = mstatusins_r[7]; // @[CSR.scala 122:75]
  wire [63:0] _mstatusval_T_2 = {mstatusval_hi_hi_hi,1'h1,mstatusval_hi_lo,mstatusval_lo_hi,mstatusval_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mstatusval_T_3 = io_rs1 | mstatusins_r; // @[CSR.scala 127:14]
  wire [63:0] _mstatusval_T_5 = _mepcval_T_2 & mstatusins_r; // @[CSR.scala 128:26]
  wire [63:0] _mstatusval_T_6 = uimmext | mstatusins_r; // @[CSR.scala 129:15]
  wire [63:0] _mstatusval_T_8 = _mepcval_T_5 & mstatusins_r; // @[CSR.scala 130:27]
  wire [63:0] _mstatusval_T_16 = sel1H[1] ? _mstatusval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_17 = sel1H[2] ? _mstatusval_T_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_18 = sel1H[3] ? _mstatusval_T_6 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_19 = sel1H[4] ? _mstatusval_T_8 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_21 = _mepcval_T_13 | _mstatusval_T_16; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_22 = _mstatusval_T_21 | _mstatusval_T_17; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_23 = _mstatusval_T_22 | _mstatusval_T_18; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_24 = _mstatusval_T_23 | _mstatusval_T_19; // @[Mux.scala 27:72]
  wire [63:0] _mstatusval_T_25 = _mstatusval_T_24 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mstatusins_T_3 = mstatusen & _mepcins_T_2; // @[CSR.scala 151:73]
  wire  miecen = csren & io_imme == 12'h304; // @[CSR.scala 153:24]
  reg [63:0] mieins_r; // @[Reg.scala 27:20]
  wire [63:0] _mieval_T = io_rs1 | mieins_r; // @[CSR.scala 159:14]
  wire [63:0] _mieval_T_2 = _mepcval_T_2 & mieins_r; // @[CSR.scala 160:26]
  wire [63:0] _mieval_T_3 = uimmext | mieins_r; // @[CSR.scala 161:15]
  wire [63:0] _mieval_T_5 = _mepcval_T_5 & mieins_r; // @[CSR.scala 162:27]
  wire [63:0] _mieval_T_13 = sel1H[1] ? _mieval_T : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_14 = sel1H[2] ? _mieval_T_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_15 = sel1H[3] ? _mieval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_16 = sel1H[4] ? _mieval_T_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_18 = _mepcval_T_13 | _mieval_T_13; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_19 = _mieval_T_18 | _mieval_T_14; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_20 = _mieval_T_19 | _mieval_T_15; // @[Mux.scala 27:72]
  wire [63:0] _mieval_T_21 = _mieval_T_20 | _mieval_T_16; // @[Mux.scala 27:72]
  wire [63:0] mieval = _mieval_T_21 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mieins_T_4 = miecen & _mtvecins_T_3; // @[CSR.scala 166:41]
  wire  mipcen = csren & io_imme == 12'h344 | intr; // @[CSR.scala 168:45]
  reg [63:0] mipins_r; // @[Reg.scala 27:20]
  wire [55:0] mipval_hi_hi = mipins_r[63:8]; // @[CSR.scala 172:15]
  wire [6:0] mipval_lo = mipins_r[6:0]; // @[CSR.scala 172:42]
  wire [63:0] _mipval_T = {mipval_hi_hi,1'h1,mipval_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mipval_T_1 = io_rs1 | mipins_r; // @[CSR.scala 177:14]
  wire [63:0] _mipval_T_3 = _mepcval_T_2 & mipins_r; // @[CSR.scala 178:26]
  wire [63:0] _mipval_T_4 = uimmext | mipins_r; // @[CSR.scala 179:15]
  wire [63:0] _mipval_T_6 = _mepcval_T_5 & mipins_r; // @[CSR.scala 180:27]
  wire [63:0] _mipval_T_14 = sel1H[1] ? _mipval_T_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_15 = sel1H[2] ? _mipval_T_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_16 = sel1H[3] ? _mipval_T_4 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_17 = sel1H[4] ? _mipval_T_6 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_19 = _mepcval_T_13 | _mipval_T_14; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_20 = _mipval_T_19 | _mipval_T_15; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_21 = _mipval_T_20 | _mipval_T_16; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_22 = _mipval_T_21 | _mipval_T_17; // @[Mux.scala 27:72]
  wire [63:0] _mipval_T_23 = _mipval_T_22 | _mepcval_T_18; // @[Mux.scala 27:72]
  wire  _mipins_T_3 = mipcen & _mepcins_T_2; // @[CSR.scala 184:42]
  wire [63:0] _io_rd_T_1 = 12'h341 == io_imme ? mepcins_r : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_rd_T_3 = 12'h342 == io_imme ? mcauseins_r : _io_rd_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_rd_T_5 = 12'h305 == io_imme ? mtvecins_r : _io_rd_T_3; // @[Mux.scala 80:57]
  wire [63:0] _io_rd_T_7 = 12'h300 == io_imme ? mstatusins_r : _io_rd_T_5; // @[Mux.scala 80:57]
  wire [63:0] _io_rd_T_9 = 12'h304 == io_imme ? mieins_r : _io_rd_T_7; // @[Mux.scala 80:57]
  wire  startTimeCnt = mieins_r[7] & mstatusval_hi_hi_lo; // @[CSR.scala 242:29]
  assign io_rd = 12'h344 == io_imme ? mipins_r : _io_rd_T_9; // @[Mux.scala 80:57]
  assign io_mtvec = mtvecins_r; // @[CSR.scala 100:22 CSR.scala 112:12]
  assign io_mepc = mepcins_r; // @[CSR.scala 59:21 CSR.scala 75:10]
  assign startTimeCnt_0 = startTimeCnt;
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      mepcins_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mepcins_T_3) begin // @[Reg.scala 28:19]
      if (_mepcval_T) begin // @[CSR.scala 60:20]
        mepcins_r <= io_pc;
      end else begin
        mepcins_r <= _mepcval_T_23;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      mcauseins_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mcauseins_T_3) begin // @[Reg.scala 28:19]
      if (intr) begin // @[CSR.scala 79:22]
        mcauseins_r <= 64'h8000000000000007;
      end else if (io_ecall) begin // @[CSR.scala 82:8]
        mcauseins_r <= 64'hb;
      end else begin
        mcauseins_r <= _mcauseval_T_22;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      mtvecins_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mtvecins_T_4) begin // @[Reg.scala 28:19]
      mtvecins_r <= mtvecval; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mstatusins_r <= 64'ha00001800; // @[Reg.scala 27:20]
    end else if (_mstatusins_T_3) begin // @[Reg.scala 28:19]
      if (_mepcval_T) begin // @[CSR.scala 117:8]
        mstatusins_r <= _mstatusval_T_1;
      end else if (io_mret) begin // @[CSR.scala 120:10]
        mstatusins_r <= _mstatusval_T_2;
      end else begin
        mstatusins_r <= _mstatusval_T_25;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      mieins_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mieins_T_4) begin // @[Reg.scala 28:19]
      mieins_r <= mieval; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mipins_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mipins_T_3) begin // @[Reg.scala 28:19]
      if (intr) begin // @[CSR.scala 170:19]
        mipins_r <= _mipval_T;
      end else begin
        mipins_r <= _mipval_T_23;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mepcins_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcauseins_r = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mtvecins_r = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatusins_r = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mieins_r = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mipins_r = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dnpcGen(
  input         io_npcSrc,
  input  [31:0] io_pc,
  input  [31:0] io_imme,
  input  [31:0] io_rd,
  output [31:0] io_dnpc
);
  wire [31:0] src1 = ~io_npcSrc ? io_rd : io_pc; // @[dnpcGen.scala 15:17]
  assign io_dnpc = io_imme + src1; // @[dnpcGen.scala 16:22]
endmodule
module memData(
  input  [63:0] io_rdata,
  output [63:0] io_rdata_ext,
  input  [2:0]  io_memReadNum
);
  wire [7:0] io_rdata_ext_lo = io_rdata[7:0]; // @[memData.scala 17:35]
  wire  io_rdata_ext_signBit = io_rdata_ext_lo[7]; // @[immeGen.scala 17:22]
  wire [55:0] io_rdata_ext_hi = io_rdata_ext_signBit ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_rdata_ext_T_1 = {io_rdata_ext_hi,io_rdata_ext_lo}; // @[Cat.scala 30:58]
  wire [15:0] io_rdata_ext_lo_1 = io_rdata[15:0]; // @[memData.scala 18:35]
  wire  io_rdata_ext_signBit_1 = io_rdata_ext_lo_1[15]; // @[immeGen.scala 17:22]
  wire [47:0] io_rdata_ext_hi_1 = io_rdata_ext_signBit_1 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_rdata_ext_T_3 = {io_rdata_ext_hi_1,io_rdata_ext_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] io_rdata_ext_lo_2 = io_rdata[31:0]; // @[memData.scala 19:35]
  wire  io_rdata_ext_signBit_2 = io_rdata_ext_lo_2[31]; // @[immeGen.scala 17:22]
  wire [31:0] io_rdata_ext_hi_2 = io_rdata_ext_signBit_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_rdata_ext_T_5 = {io_rdata_ext_hi_2,io_rdata_ext_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_rdata_ext_T_6 = {56'h0,io_rdata_ext_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_rdata_ext_T_7 = {48'h0,io_rdata_ext_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _io_rdata_ext_T_8 = {32'h0,io_rdata_ext_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_rdata_ext_T_10 = 3'h0 == io_memReadNum ? _io_rdata_ext_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_ext_T_12 = 3'h1 == io_memReadNum ? _io_rdata_ext_T_3 : _io_rdata_ext_T_10; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_ext_T_14 = 3'h2 == io_memReadNum ? _io_rdata_ext_T_5 : _io_rdata_ext_T_12; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_ext_T_16 = 3'h3 == io_memReadNum ? io_rdata : _io_rdata_ext_T_14; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_ext_T_18 = 3'h4 == io_memReadNum ? _io_rdata_ext_T_6 : _io_rdata_ext_T_16; // @[Mux.scala 80:57]
  wire [63:0] _io_rdata_ext_T_20 = 3'h5 == io_memReadNum ? _io_rdata_ext_T_7 : _io_rdata_ext_T_18; // @[Mux.scala 80:57]
  assign io_rdata_ext = 3'h6 == io_memReadNum ? _io_rdata_ext_T_8 : _io_rdata_ext_T_20; // @[Mux.scala 80:57]
endmodule
module execute(
  input          clock,
  input          reset,
  input  [1:0]   io_AluSrc1,
  input  [1:0]   io_AluSrc2,
  input  [4:0]   io_ALUCtrl,
  input          io_dnpcSrc,
  input  [1:0]   io_ResultSrc,
  input  [2:0]   io_memReadNum,
  input  [63:0]  io_dataId_imme,
  input  [63:0]  io_dataId_dOut1,
  input  [63:0]  io_dataId_dOut2,
  output [63:0]  io_dataId_dIn,
  input  [63:0]  io_dataId_rdDout,
  output [63:0]  io_dataOut_ALUResOut,
  output [63:0]  io_dataOut_wdata,
  input  [63:0]  io_dataOut_rdata,
  output         io_brTake,
  input  [31:0]  io_pc,
  input  [31:0]  io_snpc,
  output [31:0]  io_dnpc,
  input          io_CSRCtrlIf_csrrwen,
  input          io_CSRCtrlIf_csrswen,
  input          io_CSRCtrlIf_csrrsien,
  input          io_CSRCtrlIf_csrrcien,
  input          io_CSRCtrlIf_csrrcen,
  input          io_CSRCtrlIf_csrrwien,
  input          io_CSRCtrlIf_ecall,
  input          io_CSRCtrlIf_rfen,
  input          io_CSRCtrlIf_mepc2pc,
  input  [4:0]   io_uimm,
  input  [63:0]  io_aluResIn,
  input  [1:0]   io_forwardA,
  input  [1:0]   io_forwardB,
  input  [1:0]   io_forwardC,
  input  [63:0]  io_aluRes1,
  input  [63:0]  io_aluRes3,
  input          intrTimeCnt_0,
  output         startTimeCnt,
  output [191:0] dmaCtrl_0,
  input          blockDMA,
  output         block1,
  input          block23
);
  wire  ALU_clock; // @[execute.scala 97:19]
  wire  ALU_reset; // @[execute.scala 97:19]
  wire [63:0] ALU_io_srcA; // @[execute.scala 97:19]
  wire [63:0] ALU_io_srcB; // @[execute.scala 97:19]
  wire [4:0] ALU_io_ALUCtrl; // @[execute.scala 97:19]
  wire [63:0] ALU_io_ALUResult; // @[execute.scala 97:19]
  wire  ALU_block1_0; // @[execute.scala 97:19]
  wire  ALU_block23_0; // @[execute.scala 97:19]
  wire  csr_ins_clock; // @[execute.scala 104:23]
  wire  csr_ins_reset; // @[execute.scala 104:23]
  wire  csr_ins_io_csrrwen; // @[execute.scala 104:23]
  wire  csr_ins_io_csrswen; // @[execute.scala 104:23]
  wire  csr_ins_io_csrrsien; // @[execute.scala 104:23]
  wire  csr_ins_io_csrrcien; // @[execute.scala 104:23]
  wire  csr_ins_io_csrrcen; // @[execute.scala 104:23]
  wire  csr_ins_io_csrrwien; // @[execute.scala 104:23]
  wire  csr_ins_io_ecall; // @[execute.scala 104:23]
  wire [63:0] csr_ins_io_rs1; // @[execute.scala 104:23]
  wire [11:0] csr_ins_io_imme; // @[execute.scala 104:23]
  wire [63:0] csr_ins_io_pc; // @[execute.scala 104:23]
  wire [4:0] csr_ins_io_uimm; // @[execute.scala 104:23]
  wire [63:0] csr_ins_io_rd; // @[execute.scala 104:23]
  wire [63:0] csr_ins_io_mtvec; // @[execute.scala 104:23]
  wire [63:0] csr_ins_io_mepc; // @[execute.scala 104:23]
  wire  csr_ins_io_mret; // @[execute.scala 104:23]
  wire  csr_ins_intrTimeCnt_0; // @[execute.scala 104:23]
  wire  csr_ins_startTimeCnt_0; // @[execute.scala 104:23]
  wire  csr_ins_blockDMA_0; // @[execute.scala 104:23]
  wire  csr_ins_block1_0; // @[execute.scala 104:23]
  wire  csr_ins_block23_0; // @[execute.scala 104:23]
  wire  dnpcGenIns_io_npcSrc; // @[execute.scala 124:26]
  wire [31:0] dnpcGenIns_io_pc; // @[execute.scala 124:26]
  wire [31:0] dnpcGenIns_io_imme; // @[execute.scala 124:26]
  wire [31:0] dnpcGenIns_io_rd; // @[execute.scala 124:26]
  wire [31:0] dnpcGenIns_io_dnpc; // @[execute.scala 124:26]
  wire [63:0] memData_ins_io_rdata; // @[execute.scala 149:27]
  wire [63:0] memData_ins_io_rdata_ext; // @[execute.scala 149:27]
  wire [2:0] memData_ins_io_memReadNum; // @[execute.scala 149:27]
  wire [63:0] _dOut1_T_1 = 2'h2 == io_forwardA ? io_aluRes1 : io_dataId_dOut1; // @[Mux.scala 80:57]
  wire [63:0] _dinMux_T_3 = 2'h1 == io_ResultSrc ? {{32'd0}, io_snpc} : io_aluResIn; // @[Mux.scala 80:57]
  wire [63:0] dinMux = 2'h2 == io_ResultSrc ? memData_ins_io_rdata_ext : _dinMux_T_3; // @[Mux.scala 80:57]
  wire [63:0] _dOut1_T_3 = 2'h1 == io_forwardA ? dinMux : _dOut1_T_1; // @[Mux.scala 80:57]
  wire [63:0] dOut1 = 2'h3 == io_forwardA ? io_aluRes3 : _dOut1_T_3; // @[Mux.scala 80:57]
  wire [63:0] _ALUD1_T_1 = 2'h0 == io_AluSrc1 ? dOut1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _ALUD1_T_3 = 2'h1 == io_AluSrc1 ? io_dataId_imme : _ALUD1_T_1; // @[Mux.scala 80:57]
  wire [63:0] _dOut2_T_1 = 2'h2 == io_forwardB ? io_aluRes1 : io_dataId_dOut2; // @[Mux.scala 80:57]
  wire [63:0] _dOut2_T_3 = 2'h1 == io_forwardB ? dinMux : _dOut2_T_1; // @[Mux.scala 80:57]
  wire [63:0] dOut2 = 2'h3 == io_forwardB ? io_aluRes3 : _dOut2_T_3; // @[Mux.scala 80:57]
  wire [63:0] _ALUD2_T_1 = 2'h0 == io_AluSrc2 ? dOut2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _ALUD2_T_3 = 2'h1 == io_AluSrc2 ? io_dataId_imme : _ALUD2_T_1; // @[Mux.scala 80:57]
  wire [63:0] _io_dnpc_T_1 = io_CSRCtrlIf_mepc2pc ? csr_ins_io_mepc : {{32'd0}, dnpcGenIns_io_dnpc}; // @[execute.scala 135:72]
  wire [63:0] _io_dnpc_T_2 = io_CSRCtrlIf_ecall | intrTimeCnt_0 ? csr_ins_io_mtvec : _io_dnpc_T_1; // @[execute.scala 135:17]
  wire [63:0] _dmaLen_T_1 = 2'h2 == io_forwardC ? io_aluRes1 : io_dataId_rdDout; // @[Mux.scala 80:57]
  wire [63:0] _dmaLen_T_3 = 2'h1 == io_forwardC ? dinMux : _dmaLen_T_1; // @[Mux.scala 80:57]
  wire [63:0] dmaLen = 2'h3 == io_forwardC ? io_aluRes3 : _dmaLen_T_3; // @[Mux.scala 80:57]
  wire [191:0] dmaCtrl = {dmaLen,dOut2,dOut1}; // @[Cat.scala 30:58]
  ALU ALU ( // @[execute.scala 97:19]
    .clock(ALU_clock),
    .reset(ALU_reset),
    .io_srcA(ALU_io_srcA),
    .io_srcB(ALU_io_srcB),
    .io_ALUCtrl(ALU_io_ALUCtrl),
    .io_ALUResult(ALU_io_ALUResult),
    .block1_0(ALU_block1_0),
    .block23_0(ALU_block23_0)
  );
  CSR csr_ins ( // @[execute.scala 104:23]
    .clock(csr_ins_clock),
    .reset(csr_ins_reset),
    .io_csrrwen(csr_ins_io_csrrwen),
    .io_csrswen(csr_ins_io_csrswen),
    .io_csrrsien(csr_ins_io_csrrsien),
    .io_csrrcien(csr_ins_io_csrrcien),
    .io_csrrcen(csr_ins_io_csrrcen),
    .io_csrrwien(csr_ins_io_csrrwien),
    .io_ecall(csr_ins_io_ecall),
    .io_rs1(csr_ins_io_rs1),
    .io_imme(csr_ins_io_imme),
    .io_pc(csr_ins_io_pc),
    .io_uimm(csr_ins_io_uimm),
    .io_rd(csr_ins_io_rd),
    .io_mtvec(csr_ins_io_mtvec),
    .io_mepc(csr_ins_io_mepc),
    .io_mret(csr_ins_io_mret),
    .intrTimeCnt_0(csr_ins_intrTimeCnt_0),
    .startTimeCnt_0(csr_ins_startTimeCnt_0),
    .blockDMA_0(csr_ins_blockDMA_0),
    .block1_0(csr_ins_block1_0),
    .block23_0(csr_ins_block23_0)
  );
  dnpcGen dnpcGenIns ( // @[execute.scala 124:26]
    .io_npcSrc(dnpcGenIns_io_npcSrc),
    .io_pc(dnpcGenIns_io_pc),
    .io_imme(dnpcGenIns_io_imme),
    .io_rd(dnpcGenIns_io_rd),
    .io_dnpc(dnpcGenIns_io_dnpc)
  );
  memData memData_ins ( // @[execute.scala 149:27]
    .io_rdata(memData_ins_io_rdata),
    .io_rdata_ext(memData_ins_io_rdata_ext),
    .io_memReadNum(memData_ins_io_memReadNum)
  );
  assign io_dataId_dIn = 2'h2 == io_ResultSrc ? memData_ins_io_rdata_ext : _dinMux_T_3; // @[Mux.scala 80:57]
  assign io_dataOut_ALUResOut = io_CSRCtrlIf_rfen ? csr_ins_io_rd : ALU_io_ALUResult; // @[execute.scala 121:30]
  assign io_dataOut_wdata = 2'h3 == io_forwardB ? io_aluRes3 : _dOut2_T_3; // @[Mux.scala 80:57]
  assign io_brTake = ALU_io_ALUResult[0]; // @[execute.scala 137:32]
  assign io_dnpc = _io_dnpc_T_2[31:0]; // @[execute.scala 135:11]
  assign startTimeCnt = csr_ins_startTimeCnt_0;
  assign dmaCtrl_0 = dmaCtrl;
  assign block1 = ALU_block1_0;
  assign ALU_clock = clock;
  assign ALU_reset = reset;
  assign ALU_io_srcA = 2'h2 == io_AluSrc1 ? {{32'd0}, io_pc} : _ALUD1_T_3; // @[Mux.scala 80:57]
  assign ALU_io_srcB = 2'h2 == io_AluSrc2 ? {{32'd0}, io_pc} : _ALUD2_T_3; // @[Mux.scala 80:57]
  assign ALU_io_ALUCtrl = io_ALUCtrl; // @[execute.scala 100:18]
  assign ALU_block23_0 = block23;
  assign csr_ins_clock = clock;
  assign csr_ins_reset = reset;
  assign csr_ins_io_csrrwen = io_CSRCtrlIf_csrrwen; // @[execute.scala 105:22]
  assign csr_ins_io_csrswen = io_CSRCtrlIf_csrswen; // @[execute.scala 106:22]
  assign csr_ins_io_csrrsien = io_CSRCtrlIf_csrrsien; // @[execute.scala 107:23]
  assign csr_ins_io_csrrcien = io_CSRCtrlIf_csrrcien; // @[execute.scala 108:23]
  assign csr_ins_io_csrrcen = io_CSRCtrlIf_csrrcen; // @[execute.scala 109:22]
  assign csr_ins_io_csrrwien = io_CSRCtrlIf_csrrwien; // @[execute.scala 110:23]
  assign csr_ins_io_ecall = io_CSRCtrlIf_ecall; // @[execute.scala 111:20]
  assign csr_ins_io_rs1 = 2'h3 == io_forwardA ? io_aluRes3 : _dOut1_T_3; // @[Mux.scala 80:57]
  assign csr_ins_io_imme = io_dataId_imme[11:0]; // @[execute.scala 114:19]
  assign csr_ins_io_pc = {{32'd0}, io_pc}; // @[execute.scala 115:17]
  assign csr_ins_io_uimm = io_uimm; // @[execute.scala 116:19]
  assign csr_ins_io_mret = io_CSRCtrlIf_mepc2pc; // @[execute.scala 117:19]
  assign csr_ins_intrTimeCnt_0 = intrTimeCnt_0;
  assign csr_ins_blockDMA_0 = blockDMA;
  assign csr_ins_block1_0 = block1;
  assign csr_ins_block23_0 = block23;
  assign dnpcGenIns_io_npcSrc = io_dnpcSrc; // @[execute.scala 129:24]
  assign dnpcGenIns_io_pc = io_pc; // @[execute.scala 125:20]
  assign dnpcGenIns_io_imme = io_dataId_imme[31:0]; // @[execute.scala 126:22]
  assign dnpcGenIns_io_rd = dOut1[31:0]; // @[execute.scala 128:20]
  assign memData_ins_io_rdata = io_dataOut_rdata; // @[execute.scala 151:24]
  assign memData_ins_io_memReadNum = io_memReadNum; // @[execute.scala 150:29]
endmodule
module hazard(
  input        io_regEnEXMEM,
  input  [4:0] io_rdEXMEM,
  input  [4:0] io_rs1IDEX,
  input  [4:0] io_rs2IDEX,
  input        io_regEnMEMWB,
  input  [4:0] io_rdMEMWB,
  input        io_regEnWBEND,
  input  [4:0] io_rdWBEND,
  output [1:0] io_forwardA,
  output [1:0] io_forwardB,
  output [1:0] io_forwardC,
  input  [4:0] io_rs1IFID,
  input  [4:0] io_rs2IFID,
  input  [4:0] io_rdIDEX,
  input  [1:0] io_resSrc,
  output       io_loadHazard
);
  wire  _forwardAOne_T_2 = io_rs1IDEX != 5'h0; // @[hazard.scala 38:76]
  wire  forwardAOne = io_regEnEXMEM & io_rdEXMEM == io_rs1IDEX & io_rs1IDEX != 5'h0; // @[hazard.scala 38:63]
  wire  _forwardATwo_T_5 = ~io_regEnEXMEM; // @[hazard.scala 39:115]
  wire  forwardATwo = io_regEnMEMWB & io_rdMEMWB == io_rs1IDEX & _forwardAOne_T_2 & (io_rdEXMEM != io_rs1IDEX | ~
    io_regEnEXMEM); // @[hazard.scala 39:84]
  wire  forwardAThree = io_regEnWBEND & io_rdWBEND == io_rs1IDEX & _forwardAOne_T_2; // @[hazard.scala 40:66]
  wire [1:0] _io_forwardA_T = forwardAThree ? 2'h3 : 2'h0; // @[hazard.scala 41:75]
  wire [1:0] _io_forwardA_T_1 = forwardATwo ? 2'h1 : _io_forwardA_T; // @[hazard.scala 41:47]
  wire  _forwardBOne_T_2 = io_rs2IDEX != 5'h0; // @[hazard.scala 43:76]
  wire  forwardBOne = io_regEnEXMEM & io_rdEXMEM == io_rs2IDEX & io_rs2IDEX != 5'h0; // @[hazard.scala 43:63]
  wire  forwardBTwo = io_regEnMEMWB & io_rdMEMWB == io_rs2IDEX & _forwardBOne_T_2 & (io_rdEXMEM != io_rs2IDEX |
    _forwardATwo_T_5); // @[hazard.scala 44:84]
  wire  forwardBThree = io_regEnWBEND & io_rdWBEND == io_rs2IDEX & _forwardBOne_T_2; // @[hazard.scala 45:67]
  wire [1:0] _io_forwardB_T = forwardBThree ? 2'h3 : 2'h0; // @[hazard.scala 46:75]
  wire [1:0] _io_forwardB_T_1 = forwardBTwo ? 2'h1 : _io_forwardB_T; // @[hazard.scala 46:47]
  wire  _forwardCOne_T_2 = io_rdIDEX != 5'h0; // @[hazard.scala 49:76]
  wire  forwardCOne = io_regEnEXMEM & io_rdEXMEM == io_rdIDEX & io_rdIDEX != 5'h0; // @[hazard.scala 49:63]
  wire  forwardCTwo = io_regEnMEMWB & io_rdMEMWB == io_rdIDEX & _forwardCOne_T_2 & (io_rdEXMEM != io_rdIDEX |
    _forwardATwo_T_5); // @[hazard.scala 50:84]
  wire  forwardCThree = io_regEnWBEND & io_rdWBEND == io_rdIDEX & _forwardCOne_T_2; // @[hazard.scala 51:65]
  wire [1:0] _io_forwardC_T = forwardCThree ? 2'h3 : 2'h0; // @[hazard.scala 52:75]
  wire [1:0] _io_forwardC_T_1 = forwardCTwo ? 2'h1 : _io_forwardC_T; // @[hazard.scala 52:48]
  assign io_forwardA = forwardAOne ? 2'h2 : _io_forwardA_T_1; // @[hazard.scala 41:20]
  assign io_forwardB = forwardBOne ? 2'h2 : _io_forwardB_T_1; // @[hazard.scala 46:21]
  assign io_forwardC = forwardCOne ? 2'h2 : _io_forwardC_T_1; // @[hazard.scala 52:21]
  assign io_loadHazard = (io_rs1IFID == io_rdIDEX | io_rs2IFID == io_rdIDEX) & io_resSrc == 2'h2; // @[hazard.scala 57:74]
endmodule
module preCell(
  input         clock,
  input         reset,
  input         io_cen,
  input         io_jump,
  input  [31:0] io_dnpcIn,
  output [31:0] io_dnpcOut,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _dnpcReg_T = io_cen & io_jump; // @[preCell.scala 16:48]
  reg [31:0] dnpcReg; // @[Reg.scala 27:20]
  wire  takenV = dnpcReg == io_dnpcIn; // @[preCell.scala 21:24]
  wire [1:0] sntMux = takenV ? 2'h1 : 2'h0; // @[preCell.scala 22:19]
  wire [1:0] ntMux = takenV ? 2'h2 : 2'h0; // @[preCell.scala 23:18]
  wire [1:0] tMux = takenV ? 2'h3 : 2'h1; // @[preCell.scala 24:17]
  reg [1:0] stateWire_r; // @[Reg.scala 27:20]
  wire [1:0] _stateWire_T_1 = 2'h1 == stateWire_r ? ntMux : sntMux; // @[Mux.scala 80:57]
  assign io_dnpcOut = dnpcReg; // @[preCell.scala 42:14]
  assign io_valid = stateWire_r == 2'h2 | stateWire_r == 2'h3; // @[preCell.scala 43:35]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      dnpcReg <= 32'h0; // @[Reg.scala 27:20]
    end else if (_dnpcReg_T) begin // @[Reg.scala 28:19]
      dnpcReg <= io_dnpcIn; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      stateWire_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (io_cen) begin // @[Reg.scala 28:19]
      if (2'h3 == stateWire_r) begin // @[Mux.scala 80:57]
        if (takenV) begin // @[preCell.scala 25:18]
          stateWire_r <= 2'h3;
        end else begin
          stateWire_r <= 2'h2;
        end
      end else if (2'h2 == stateWire_r) begin // @[Mux.scala 80:57]
        stateWire_r <= tMux;
      end else begin
        stateWire_r <= _stateWire_T_1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dnpcReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stateWire_r = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module preBranch(
  input         clock,
  input         reset,
  input         io_exjump,
  input  [31:0] io_ifpc,
  input  [31:0] io_expc,
  input  [31:0] io_exdpc,
  output [31:0] io_ifdnpc,
  output        io_ifjump,
  input         block1_0,
  input         block23_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  precelList_0_clock; // @[preBranch.scala 29:45]
  wire  precelList_0_reset; // @[preBranch.scala 29:45]
  wire  precelList_0_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_0_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_0_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_0_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_0_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_1_clock; // @[preBranch.scala 29:45]
  wire  precelList_1_reset; // @[preBranch.scala 29:45]
  wire  precelList_1_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_1_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_1_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_1_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_1_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_2_clock; // @[preBranch.scala 29:45]
  wire  precelList_2_reset; // @[preBranch.scala 29:45]
  wire  precelList_2_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_2_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_2_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_2_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_2_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_3_clock; // @[preBranch.scala 29:45]
  wire  precelList_3_reset; // @[preBranch.scala 29:45]
  wire  precelList_3_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_3_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_3_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_3_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_3_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_4_clock; // @[preBranch.scala 29:45]
  wire  precelList_4_reset; // @[preBranch.scala 29:45]
  wire  precelList_4_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_4_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_4_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_4_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_4_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_5_clock; // @[preBranch.scala 29:45]
  wire  precelList_5_reset; // @[preBranch.scala 29:45]
  wire  precelList_5_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_5_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_5_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_5_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_5_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_6_clock; // @[preBranch.scala 29:45]
  wire  precelList_6_reset; // @[preBranch.scala 29:45]
  wire  precelList_6_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_6_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_6_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_6_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_6_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_7_clock; // @[preBranch.scala 29:45]
  wire  precelList_7_reset; // @[preBranch.scala 29:45]
  wire  precelList_7_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_7_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_7_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_7_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_7_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_8_clock; // @[preBranch.scala 29:45]
  wire  precelList_8_reset; // @[preBranch.scala 29:45]
  wire  precelList_8_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_8_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_8_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_8_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_8_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_9_clock; // @[preBranch.scala 29:45]
  wire  precelList_9_reset; // @[preBranch.scala 29:45]
  wire  precelList_9_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_9_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_9_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_9_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_9_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_10_clock; // @[preBranch.scala 29:45]
  wire  precelList_10_reset; // @[preBranch.scala 29:45]
  wire  precelList_10_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_10_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_10_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_10_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_10_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_11_clock; // @[preBranch.scala 29:45]
  wire  precelList_11_reset; // @[preBranch.scala 29:45]
  wire  precelList_11_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_11_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_11_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_11_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_11_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_12_clock; // @[preBranch.scala 29:45]
  wire  precelList_12_reset; // @[preBranch.scala 29:45]
  wire  precelList_12_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_12_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_12_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_12_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_12_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_13_clock; // @[preBranch.scala 29:45]
  wire  precelList_13_reset; // @[preBranch.scala 29:45]
  wire  precelList_13_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_13_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_13_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_13_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_13_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_14_clock; // @[preBranch.scala 29:45]
  wire  precelList_14_reset; // @[preBranch.scala 29:45]
  wire  precelList_14_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_14_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_14_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_14_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_14_io_valid; // @[preBranch.scala 29:45]
  wire  precelList_15_clock; // @[preBranch.scala 29:45]
  wire  precelList_15_reset; // @[preBranch.scala 29:45]
  wire  precelList_15_io_cen; // @[preBranch.scala 29:45]
  wire  precelList_15_io_jump; // @[preBranch.scala 29:45]
  wire [31:0] precelList_15_io_dnpcIn; // @[preBranch.scala 29:45]
  wire [31:0] precelList_15_io_dnpcOut; // @[preBranch.scala 29:45]
  wire  precelList_15_io_valid; // @[preBranch.scala 29:45]
  wire  block = block1_0 | block23_0; // @[preBranch.scala 26:33]
  reg [31:0] pcList_0_r; // @[Reg.scala 27:20]
  reg  vList_0_r; // @[Reg.scala 27:20]
  wire  hitList_0 = io_expc == pcList_0_r & vList_0_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_1_r; // @[Reg.scala 27:20]
  reg  vList_1_r; // @[Reg.scala 27:20]
  wire  hitList_1 = io_expc == pcList_1_r & vList_1_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_2_r; // @[Reg.scala 27:20]
  reg  vList_2_r; // @[Reg.scala 27:20]
  wire  hitList_2 = io_expc == pcList_2_r & vList_2_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_3_r; // @[Reg.scala 27:20]
  reg  vList_3_r; // @[Reg.scala 27:20]
  wire  hitList_3 = io_expc == pcList_3_r & vList_3_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_4_r; // @[Reg.scala 27:20]
  reg  vList_4_r; // @[Reg.scala 27:20]
  wire  hitList_4 = io_expc == pcList_4_r & vList_4_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_5_r; // @[Reg.scala 27:20]
  reg  vList_5_r; // @[Reg.scala 27:20]
  wire  hitList_5 = io_expc == pcList_5_r & vList_5_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_6_r; // @[Reg.scala 27:20]
  reg  vList_6_r; // @[Reg.scala 27:20]
  wire  hitList_6 = io_expc == pcList_6_r & vList_6_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_7_r; // @[Reg.scala 27:20]
  reg  vList_7_r; // @[Reg.scala 27:20]
  wire  hitList_7 = io_expc == pcList_7_r & vList_7_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_8_r; // @[Reg.scala 27:20]
  reg  vList_8_r; // @[Reg.scala 27:20]
  wire  hitList_8 = io_expc == pcList_8_r & vList_8_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_9_r; // @[Reg.scala 27:20]
  reg  vList_9_r; // @[Reg.scala 27:20]
  wire  hitList_9 = io_expc == pcList_9_r & vList_9_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_10_r; // @[Reg.scala 27:20]
  reg  vList_10_r; // @[Reg.scala 27:20]
  wire  hitList_10 = io_expc == pcList_10_r & vList_10_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_11_r; // @[Reg.scala 27:20]
  reg  vList_11_r; // @[Reg.scala 27:20]
  wire  hitList_11 = io_expc == pcList_11_r & vList_11_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_12_r; // @[Reg.scala 27:20]
  reg  vList_12_r; // @[Reg.scala 27:20]
  wire  hitList_12 = io_expc == pcList_12_r & vList_12_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_13_r; // @[Reg.scala 27:20]
  reg  vList_13_r; // @[Reg.scala 27:20]
  wire  hitList_13 = io_expc == pcList_13_r & vList_13_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_14_r; // @[Reg.scala 27:20]
  reg  vList_14_r; // @[Reg.scala 27:20]
  wire  hitList_14 = io_expc == pcList_14_r & vList_14_r; // @[preBranch.scala 35:41]
  reg [31:0] pcList_15_r; // @[Reg.scala 27:20]
  reg  vList_15_r; // @[Reg.scala 27:20]
  wire  hitList_15 = io_expc == pcList_15_r & vList_15_r; // @[preBranch.scala 35:41]
  wire  hit = hitList_0 | hitList_1 | hitList_2 | hitList_3 | hitList_4 | hitList_5 | hitList_6 | hitList_7 | hitList_8
     | hitList_9 | hitList_10 | hitList_11 | hitList_12 | hitList_13 | hitList_14 | hitList_15; // @[preBranch.scala 37:51]
  reg [3:0] cnt_r; // @[Reg.scala 27:20]
  wire [3:0] _cnt_T_1 = cnt_r + 4'h1; // @[preBranch.scala 40:25]
  wire  _cnt_T_4 = ~block; // @[preBranch.scala 40:61]
  wire  _cnt_T_5 = ~hit & io_exjump & ~block; // @[preBranch.scala 40:58]
  wire  _precelList_0_io_cen_T = cnt_r == 4'h0; // @[preBranch.scala 46:62]
  wire  _vList_0_T_5 = ~hitList_0 & io_exjump & _precelList_0_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_1 = _vList_0_T_5 | vList_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_1_io_cen_T = cnt_r == 4'h1; // @[preBranch.scala 46:62]
  wire  _vList_1_T_5 = ~hitList_1 & io_exjump & _precelList_1_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_3 = _vList_1_T_5 | vList_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_2_io_cen_T = cnt_r == 4'h2; // @[preBranch.scala 46:62]
  wire  _vList_2_T_5 = ~hitList_2 & io_exjump & _precelList_2_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_5 = _vList_2_T_5 | vList_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_3_io_cen_T = cnt_r == 4'h3; // @[preBranch.scala 46:62]
  wire  _vList_3_T_5 = ~hitList_3 & io_exjump & _precelList_3_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_7 = _vList_3_T_5 | vList_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_4_io_cen_T = cnt_r == 4'h4; // @[preBranch.scala 46:62]
  wire  _vList_4_T_5 = ~hitList_4 & io_exjump & _precelList_4_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_9 = _vList_4_T_5 | vList_4_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_5_io_cen_T = cnt_r == 4'h5; // @[preBranch.scala 46:62]
  wire  _vList_5_T_5 = ~hitList_5 & io_exjump & _precelList_5_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_11 = _vList_5_T_5 | vList_5_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_6_io_cen_T = cnt_r == 4'h6; // @[preBranch.scala 46:62]
  wire  _vList_6_T_5 = ~hitList_6 & io_exjump & _precelList_6_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_13 = _vList_6_T_5 | vList_6_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_7_io_cen_T = cnt_r == 4'h7; // @[preBranch.scala 46:62]
  wire  _vList_7_T_5 = ~hitList_7 & io_exjump & _precelList_7_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_15 = _vList_7_T_5 | vList_7_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_8_io_cen_T = cnt_r == 4'h8; // @[preBranch.scala 46:62]
  wire  _vList_8_T_5 = ~hitList_8 & io_exjump & _precelList_8_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_17 = _vList_8_T_5 | vList_8_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_9_io_cen_T = cnt_r == 4'h9; // @[preBranch.scala 46:62]
  wire  _vList_9_T_5 = ~hitList_9 & io_exjump & _precelList_9_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_19 = _vList_9_T_5 | vList_9_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_10_io_cen_T = cnt_r == 4'ha; // @[preBranch.scala 46:62]
  wire  _vList_10_T_5 = ~hitList_10 & io_exjump & _precelList_10_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_21 = _vList_10_T_5 | vList_10_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_11_io_cen_T = cnt_r == 4'hb; // @[preBranch.scala 46:62]
  wire  _vList_11_T_5 = ~hitList_11 & io_exjump & _precelList_11_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_23 = _vList_11_T_5 | vList_11_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_12_io_cen_T = cnt_r == 4'hc; // @[preBranch.scala 46:62]
  wire  _vList_12_T_5 = ~hitList_12 & io_exjump & _precelList_12_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_25 = _vList_12_T_5 | vList_12_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_13_io_cen_T = cnt_r == 4'hd; // @[preBranch.scala 46:62]
  wire  _vList_13_T_5 = ~hitList_13 & io_exjump & _precelList_13_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_27 = _vList_13_T_5 | vList_13_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_14_io_cen_T = cnt_r == 4'he; // @[preBranch.scala 46:62]
  wire  _vList_14_T_5 = ~hitList_14 & io_exjump & _precelList_14_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_29 = _vList_14_T_5 | vList_14_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _precelList_15_io_cen_T = cnt_r == 4'hf; // @[preBranch.scala 46:62]
  wire  _vList_15_T_5 = ~hitList_15 & io_exjump & _precelList_15_io_cen_T & _cnt_T_4; // @[preBranch.scala 48:82]
  wire  _GEN_31 = _vList_15_T_5 | vList_15_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  hitIfList_0 = io_ifpc == pcList_0_r & vList_0_r; // @[preBranch.scala 57:43]
  wire  hitIfList_1 = io_ifpc == pcList_1_r & vList_1_r; // @[preBranch.scala 57:43]
  wire  hitIfList_2 = io_ifpc == pcList_2_r & vList_2_r; // @[preBranch.scala 57:43]
  wire  hitIfList_3 = io_ifpc == pcList_3_r & vList_3_r; // @[preBranch.scala 57:43]
  wire  hitIfList_4 = io_ifpc == pcList_4_r & vList_4_r; // @[preBranch.scala 57:43]
  wire  hitIfList_5 = io_ifpc == pcList_5_r & vList_5_r; // @[preBranch.scala 57:43]
  wire  hitIfList_6 = io_ifpc == pcList_6_r & vList_6_r; // @[preBranch.scala 57:43]
  wire  hitIfList_7 = io_ifpc == pcList_7_r & vList_7_r; // @[preBranch.scala 57:43]
  wire  hitIfList_8 = io_ifpc == pcList_8_r & vList_8_r; // @[preBranch.scala 57:43]
  wire  hitIfList_9 = io_ifpc == pcList_9_r & vList_9_r; // @[preBranch.scala 57:43]
  wire  hitIfList_10 = io_ifpc == pcList_10_r & vList_10_r; // @[preBranch.scala 57:43]
  wire  hitIfList_11 = io_ifpc == pcList_11_r & vList_11_r; // @[preBranch.scala 57:43]
  wire  hitIfList_12 = io_ifpc == pcList_12_r & vList_12_r; // @[preBranch.scala 57:43]
  wire  hitIfList_13 = io_ifpc == pcList_13_r & vList_13_r; // @[preBranch.scala 57:43]
  wire  hitIfList_14 = io_ifpc == pcList_14_r & vList_14_r; // @[preBranch.scala 57:43]
  wire  hitIfList_15 = io_ifpc == pcList_15_r & vList_15_r; // @[preBranch.scala 57:43]
  wire  hitif = hitIfList_0 | hitIfList_1 | hitIfList_2 | hitIfList_3 | hitIfList_4 | hitIfList_5 | hitIfList_6 |
    hitIfList_7 | hitIfList_8 | hitIfList_9 | hitIfList_10 | hitIfList_11 | hitIfList_12 | hitIfList_13 | hitIfList_14
     | hitIfList_15; // @[preBranch.scala 60:55]
  wire  _io_ifjump_T = ~hitif; // @[preBranch.scala 66:5]
  wire  _io_ifjump_T_16 = hitIfList_15 & precelList_15_io_valid; // @[Mux.scala 27:72]
  wire  _io_ifjump_T_31 = hitIfList_0 & precelList_0_io_valid | hitIfList_1 & precelList_1_io_valid | hitIfList_2 &
    precelList_2_io_valid | hitIfList_3 & precelList_3_io_valid | hitIfList_4 & precelList_4_io_valid | hitIfList_5 &
    precelList_5_io_valid | hitIfList_6 & precelList_6_io_valid | hitIfList_7 & precelList_7_io_valid | hitIfList_8 &
    precelList_8_io_valid | hitIfList_9 & precelList_9_io_valid | hitIfList_10 & precelList_10_io_valid | hitIfList_11
     & precelList_11_io_valid | hitIfList_12 & precelList_12_io_valid | hitIfList_13 & precelList_13_io_valid |
    hitIfList_14 & precelList_14_io_valid | _io_ifjump_T_16; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_1 = hitIfList_0 ? precelList_0_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_2 = hitIfList_1 ? precelList_1_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_3 = hitIfList_2 ? precelList_2_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_4 = hitIfList_3 ? precelList_3_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_5 = hitIfList_4 ? precelList_4_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_6 = hitIfList_5 ? precelList_5_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_7 = hitIfList_6 ? precelList_6_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_8 = hitIfList_7 ? precelList_7_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_9 = hitIfList_8 ? precelList_8_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_10 = hitIfList_9 ? precelList_9_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_11 = hitIfList_10 ? precelList_10_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_12 = hitIfList_11 ? precelList_11_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_13 = hitIfList_12 ? precelList_12_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_14 = hitIfList_13 ? precelList_13_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_15 = hitIfList_14 ? precelList_14_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_16 = hitIfList_15 ? precelList_15_io_dnpcOut : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_17 = _io_ifdnpc_T_1 | _io_ifdnpc_T_2; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_18 = _io_ifdnpc_T_17 | _io_ifdnpc_T_3; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_19 = _io_ifdnpc_T_18 | _io_ifdnpc_T_4; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_20 = _io_ifdnpc_T_19 | _io_ifdnpc_T_5; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_21 = _io_ifdnpc_T_20 | _io_ifdnpc_T_6; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_22 = _io_ifdnpc_T_21 | _io_ifdnpc_T_7; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_23 = _io_ifdnpc_T_22 | _io_ifdnpc_T_8; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_24 = _io_ifdnpc_T_23 | _io_ifdnpc_T_9; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_25 = _io_ifdnpc_T_24 | _io_ifdnpc_T_10; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_26 = _io_ifdnpc_T_25 | _io_ifdnpc_T_11; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_27 = _io_ifdnpc_T_26 | _io_ifdnpc_T_12; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_28 = _io_ifdnpc_T_27 | _io_ifdnpc_T_13; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_29 = _io_ifdnpc_T_28 | _io_ifdnpc_T_14; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_30 = _io_ifdnpc_T_29 | _io_ifdnpc_T_15; // @[Mux.scala 27:72]
  wire [31:0] _io_ifdnpc_T_31 = _io_ifdnpc_T_30 | _io_ifdnpc_T_16; // @[Mux.scala 27:72]
  preCell precelList_0 ( // @[preBranch.scala 29:45]
    .clock(precelList_0_clock),
    .reset(precelList_0_reset),
    .io_cen(precelList_0_io_cen),
    .io_jump(precelList_0_io_jump),
    .io_dnpcIn(precelList_0_io_dnpcIn),
    .io_dnpcOut(precelList_0_io_dnpcOut),
    .io_valid(precelList_0_io_valid)
  );
  preCell precelList_1 ( // @[preBranch.scala 29:45]
    .clock(precelList_1_clock),
    .reset(precelList_1_reset),
    .io_cen(precelList_1_io_cen),
    .io_jump(precelList_1_io_jump),
    .io_dnpcIn(precelList_1_io_dnpcIn),
    .io_dnpcOut(precelList_1_io_dnpcOut),
    .io_valid(precelList_1_io_valid)
  );
  preCell precelList_2 ( // @[preBranch.scala 29:45]
    .clock(precelList_2_clock),
    .reset(precelList_2_reset),
    .io_cen(precelList_2_io_cen),
    .io_jump(precelList_2_io_jump),
    .io_dnpcIn(precelList_2_io_dnpcIn),
    .io_dnpcOut(precelList_2_io_dnpcOut),
    .io_valid(precelList_2_io_valid)
  );
  preCell precelList_3 ( // @[preBranch.scala 29:45]
    .clock(precelList_3_clock),
    .reset(precelList_3_reset),
    .io_cen(precelList_3_io_cen),
    .io_jump(precelList_3_io_jump),
    .io_dnpcIn(precelList_3_io_dnpcIn),
    .io_dnpcOut(precelList_3_io_dnpcOut),
    .io_valid(precelList_3_io_valid)
  );
  preCell precelList_4 ( // @[preBranch.scala 29:45]
    .clock(precelList_4_clock),
    .reset(precelList_4_reset),
    .io_cen(precelList_4_io_cen),
    .io_jump(precelList_4_io_jump),
    .io_dnpcIn(precelList_4_io_dnpcIn),
    .io_dnpcOut(precelList_4_io_dnpcOut),
    .io_valid(precelList_4_io_valid)
  );
  preCell precelList_5 ( // @[preBranch.scala 29:45]
    .clock(precelList_5_clock),
    .reset(precelList_5_reset),
    .io_cen(precelList_5_io_cen),
    .io_jump(precelList_5_io_jump),
    .io_dnpcIn(precelList_5_io_dnpcIn),
    .io_dnpcOut(precelList_5_io_dnpcOut),
    .io_valid(precelList_5_io_valid)
  );
  preCell precelList_6 ( // @[preBranch.scala 29:45]
    .clock(precelList_6_clock),
    .reset(precelList_6_reset),
    .io_cen(precelList_6_io_cen),
    .io_jump(precelList_6_io_jump),
    .io_dnpcIn(precelList_6_io_dnpcIn),
    .io_dnpcOut(precelList_6_io_dnpcOut),
    .io_valid(precelList_6_io_valid)
  );
  preCell precelList_7 ( // @[preBranch.scala 29:45]
    .clock(precelList_7_clock),
    .reset(precelList_7_reset),
    .io_cen(precelList_7_io_cen),
    .io_jump(precelList_7_io_jump),
    .io_dnpcIn(precelList_7_io_dnpcIn),
    .io_dnpcOut(precelList_7_io_dnpcOut),
    .io_valid(precelList_7_io_valid)
  );
  preCell precelList_8 ( // @[preBranch.scala 29:45]
    .clock(precelList_8_clock),
    .reset(precelList_8_reset),
    .io_cen(precelList_8_io_cen),
    .io_jump(precelList_8_io_jump),
    .io_dnpcIn(precelList_8_io_dnpcIn),
    .io_dnpcOut(precelList_8_io_dnpcOut),
    .io_valid(precelList_8_io_valid)
  );
  preCell precelList_9 ( // @[preBranch.scala 29:45]
    .clock(precelList_9_clock),
    .reset(precelList_9_reset),
    .io_cen(precelList_9_io_cen),
    .io_jump(precelList_9_io_jump),
    .io_dnpcIn(precelList_9_io_dnpcIn),
    .io_dnpcOut(precelList_9_io_dnpcOut),
    .io_valid(precelList_9_io_valid)
  );
  preCell precelList_10 ( // @[preBranch.scala 29:45]
    .clock(precelList_10_clock),
    .reset(precelList_10_reset),
    .io_cen(precelList_10_io_cen),
    .io_jump(precelList_10_io_jump),
    .io_dnpcIn(precelList_10_io_dnpcIn),
    .io_dnpcOut(precelList_10_io_dnpcOut),
    .io_valid(precelList_10_io_valid)
  );
  preCell precelList_11 ( // @[preBranch.scala 29:45]
    .clock(precelList_11_clock),
    .reset(precelList_11_reset),
    .io_cen(precelList_11_io_cen),
    .io_jump(precelList_11_io_jump),
    .io_dnpcIn(precelList_11_io_dnpcIn),
    .io_dnpcOut(precelList_11_io_dnpcOut),
    .io_valid(precelList_11_io_valid)
  );
  preCell precelList_12 ( // @[preBranch.scala 29:45]
    .clock(precelList_12_clock),
    .reset(precelList_12_reset),
    .io_cen(precelList_12_io_cen),
    .io_jump(precelList_12_io_jump),
    .io_dnpcIn(precelList_12_io_dnpcIn),
    .io_dnpcOut(precelList_12_io_dnpcOut),
    .io_valid(precelList_12_io_valid)
  );
  preCell precelList_13 ( // @[preBranch.scala 29:45]
    .clock(precelList_13_clock),
    .reset(precelList_13_reset),
    .io_cen(precelList_13_io_cen),
    .io_jump(precelList_13_io_jump),
    .io_dnpcIn(precelList_13_io_dnpcIn),
    .io_dnpcOut(precelList_13_io_dnpcOut),
    .io_valid(precelList_13_io_valid)
  );
  preCell precelList_14 ( // @[preBranch.scala 29:45]
    .clock(precelList_14_clock),
    .reset(precelList_14_reset),
    .io_cen(precelList_14_io_cen),
    .io_jump(precelList_14_io_jump),
    .io_dnpcIn(precelList_14_io_dnpcIn),
    .io_dnpcOut(precelList_14_io_dnpcOut),
    .io_valid(precelList_14_io_valid)
  );
  preCell precelList_15 ( // @[preBranch.scala 29:45]
    .clock(precelList_15_clock),
    .reset(precelList_15_reset),
    .io_cen(precelList_15_io_cen),
    .io_jump(precelList_15_io_jump),
    .io_dnpcIn(precelList_15_io_dnpcIn),
    .io_dnpcOut(precelList_15_io_dnpcOut),
    .io_valid(precelList_15_io_valid)
  );
  assign io_ifdnpc = _io_ifjump_T ? 32'h0 : _io_ifdnpc_T_31; // @[preBranch.scala 77:19]
  assign io_ifjump = _io_ifjump_T ? 1'h0 : _io_ifjump_T_31; // @[preBranch.scala 65:18]
  assign precelList_0_clock = clock;
  assign precelList_0_reset = reset;
  assign precelList_0_io_cen = (hitList_0 | io_exjump & cnt_r == 4'h0) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_0_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_0_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_1_clock = clock;
  assign precelList_1_reset = reset;
  assign precelList_1_io_cen = (hitList_1 | io_exjump & cnt_r == 4'h1) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_1_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_1_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_2_clock = clock;
  assign precelList_2_reset = reset;
  assign precelList_2_io_cen = (hitList_2 | io_exjump & cnt_r == 4'h2) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_2_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_2_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_3_clock = clock;
  assign precelList_3_reset = reset;
  assign precelList_3_io_cen = (hitList_3 | io_exjump & cnt_r == 4'h3) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_3_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_3_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_4_clock = clock;
  assign precelList_4_reset = reset;
  assign precelList_4_io_cen = (hitList_4 | io_exjump & cnt_r == 4'h4) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_4_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_4_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_5_clock = clock;
  assign precelList_5_reset = reset;
  assign precelList_5_io_cen = (hitList_5 | io_exjump & cnt_r == 4'h5) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_5_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_5_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_6_clock = clock;
  assign precelList_6_reset = reset;
  assign precelList_6_io_cen = (hitList_6 | io_exjump & cnt_r == 4'h6) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_6_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_6_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_7_clock = clock;
  assign precelList_7_reset = reset;
  assign precelList_7_io_cen = (hitList_7 | io_exjump & cnt_r == 4'h7) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_7_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_7_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_8_clock = clock;
  assign precelList_8_reset = reset;
  assign precelList_8_io_cen = (hitList_8 | io_exjump & cnt_r == 4'h8) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_8_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_8_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_9_clock = clock;
  assign precelList_9_reset = reset;
  assign precelList_9_io_cen = (hitList_9 | io_exjump & cnt_r == 4'h9) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_9_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_9_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_10_clock = clock;
  assign precelList_10_reset = reset;
  assign precelList_10_io_cen = (hitList_10 | io_exjump & cnt_r == 4'ha) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_10_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_10_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_11_clock = clock;
  assign precelList_11_reset = reset;
  assign precelList_11_io_cen = (hitList_11 | io_exjump & cnt_r == 4'hb) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_11_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_11_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_12_clock = clock;
  assign precelList_12_reset = reset;
  assign precelList_12_io_cen = (hitList_12 | io_exjump & cnt_r == 4'hc) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_12_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_12_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_13_clock = clock;
  assign precelList_13_reset = reset;
  assign precelList_13_io_cen = (hitList_13 | io_exjump & cnt_r == 4'hd) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_13_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_13_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_14_clock = clock;
  assign precelList_14_reset = reset;
  assign precelList_14_io_cen = (hitList_14 | io_exjump & cnt_r == 4'he) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_14_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_14_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  assign precelList_15_clock = clock;
  assign precelList_15_reset = reset;
  assign precelList_15_io_cen = (hitList_15 | io_exjump & cnt_r == 4'hf) & _cnt_T_4; // @[preBranch.scala 46:72]
  assign precelList_15_io_jump = io_exjump; // @[preBranch.scala 44:27]
  assign precelList_15_io_dnpcIn = io_exdpc; // @[preBranch.scala 45:29]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      pcList_0_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_0_T_5) begin // @[Reg.scala 28:19]
      pcList_0_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_0_r <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_1_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_1_T_5) begin // @[Reg.scala 28:19]
      pcList_1_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_1_r <= _GEN_3;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_2_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_2_T_5) begin // @[Reg.scala 28:19]
      pcList_2_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_2_r <= _GEN_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_3_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_3_T_5) begin // @[Reg.scala 28:19]
      pcList_3_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_3_r <= _GEN_7;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_4_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_4_T_5) begin // @[Reg.scala 28:19]
      pcList_4_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_4_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_4_r <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_5_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_5_T_5) begin // @[Reg.scala 28:19]
      pcList_5_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_5_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_5_r <= _GEN_11;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_6_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_6_T_5) begin // @[Reg.scala 28:19]
      pcList_6_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_6_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_6_r <= _GEN_13;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_7_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_7_T_5) begin // @[Reg.scala 28:19]
      pcList_7_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_7_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_7_r <= _GEN_15;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_8_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_8_T_5) begin // @[Reg.scala 28:19]
      pcList_8_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_8_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_8_r <= _GEN_17;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_9_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_9_T_5) begin // @[Reg.scala 28:19]
      pcList_9_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_9_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_9_r <= _GEN_19;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_10_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_10_T_5) begin // @[Reg.scala 28:19]
      pcList_10_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_10_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_10_r <= _GEN_21;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_11_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_11_T_5) begin // @[Reg.scala 28:19]
      pcList_11_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_11_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_11_r <= _GEN_23;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_12_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_12_T_5) begin // @[Reg.scala 28:19]
      pcList_12_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_12_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_12_r <= _GEN_25;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_13_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_13_T_5) begin // @[Reg.scala 28:19]
      pcList_13_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_13_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_13_r <= _GEN_27;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_14_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_14_T_5) begin // @[Reg.scala 28:19]
      pcList_14_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_14_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_14_r <= _GEN_29;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcList_15_r <= 32'h0; // @[Reg.scala 27:20]
    end else if (_vList_15_T_5) begin // @[Reg.scala 28:19]
      pcList_15_r <= io_expc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vList_15_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vList_15_r <= _GEN_31;
    end
    if (reset) begin // @[Reg.scala 27:20]
      cnt_r <= 4'h0; // @[Reg.scala 27:20]
    end else if (_cnt_T_5) begin // @[Reg.scala 28:19]
      cnt_r <= _cnt_T_1; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcList_0_r = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  vList_0_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pcList_1_r = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  vList_1_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pcList_2_r = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  vList_2_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pcList_3_r = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  vList_3_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pcList_4_r = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  vList_4_r = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pcList_5_r = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  vList_5_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pcList_6_r = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  vList_6_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pcList_7_r = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  vList_7_r = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pcList_8_r = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  vList_8_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pcList_9_r = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  vList_9_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pcList_10_r = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  vList_10_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pcList_11_r = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  vList_11_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  pcList_12_r = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  vList_12_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pcList_13_r = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  vList_13_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  pcList_14_r = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  vList_14_r = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pcList_15_r = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  vList_15_r = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cnt_r = _RAND_32[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module memVGen(
  input  [31:0] io_inst,
  output        io_valid
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memVGen.scala 20:45]
  wire  _T_1 = 32'h3023 == _T; // @[memVGen.scala 20:45]
  wire  _T_3 = 32'h23 == _T; // @[memVGen.scala 20:45]
  wire  _T_5 = 32'h2023 == _T; // @[memVGen.scala 20:45]
  wire  _T_7 = 32'h1023 == _T; // @[memVGen.scala 20:45]
  wire  _T_9 = 32'h3003 == _T; // @[memVGen.scala 26:27]
  wire  _T_11 = 32'h4003 == _T; // @[memVGen.scala 27:27]
  wire  _T_13 = 32'h1003 == _T; // @[memVGen.scala 28:27]
  wire  _T_15 = 32'h2003 == _T; // @[memVGen.scala 29:27]
  wire  _T_19 = 32'h5003 == _T; // @[memVGen.scala 31:27]
  wire  _T_21 = 32'h3 == _T; // @[memVGen.scala 32:27]
  wire  _T_23 = 32'h6003 == _T; // @[memVGen.scala 33:27]
  assign io_valid = _T_1 | (_T_3 | (_T_5 | (_T_7 | (_T_9 | (_T_11 | (_T_13 | (_T_15 | (_T_9 | (_T_19 | (_T_21 | _T_23)))
    ))))))); // @[Mux.scala 98:16]
endmodule
module ALUCtrl(
  input  [31:0] io_inst,
  output [4:0]  io_ALUCtrl
);
  wire [31:0] _T = io_inst & 32'h707f; // @[ALUCtrl.scala 74:49]
  wire  _T_1 = 32'h3023 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_3 = 32'h23 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_5 = 32'h2023 == _T; // @[ALUCtrl.scala 74:49]
  wire  _T_7 = 32'h1023 == _T; // @[ALUCtrl.scala 74:49]
  wire [31:0] _T_8 = io_inst & 32'h7f; // @[ALUCtrl.scala 79:31]
  wire  _T_9 = 32'h17 == _T_8; // @[ALUCtrl.scala 79:31]
  wire  _T_11 = 32'h37 == _T_8; // @[ALUCtrl.scala 80:31]
  wire  _T_13 = 32'h13 == _T; // @[ALUCtrl.scala 81:31]
  wire  _T_15 = 32'h67 == _T; // @[ALUCtrl.scala 82:31]
  wire  _T_17 = 32'h3003 == _T; // @[ALUCtrl.scala 83:31]
  wire  _T_19 = 32'h4003 == _T; // @[ALUCtrl.scala 84:31]
  wire  _T_21 = 32'h3013 == _T; // @[ALUCtrl.scala 85:31]
  wire [31:0] _T_22 = io_inst & 32'hfe00707f; // @[ALUCtrl.scala 86:31]
  wire  _T_23 = 32'h501b == _T_22; // @[ALUCtrl.scala 86:31]
  wire [31:0] _T_24 = io_inst & 32'hfc00707f; // @[ALUCtrl.scala 87:31]
  wire  _T_25 = 32'h1013 == _T_24; // @[ALUCtrl.scala 87:31]
  wire  _T_27 = 32'h7013 == _T; // @[ALUCtrl.scala 88:31]
  wire  _T_29 = 32'h4013 == _T; // @[ALUCtrl.scala 89:31]
  wire  _T_31 = 32'h1b == _T; // @[ALUCtrl.scala 90:31]
  wire  _T_33 = 32'h5013 == _T_24; // @[ALUCtrl.scala 91:31]
  wire  _T_35 = 32'h101b == _T_22; // @[ALUCtrl.scala 92:31]
  wire  _T_37 = 32'h4000501b == _T_22; // @[ALUCtrl.scala 93:31]
  wire  _T_39 = 32'h40005013 == _T_24; // @[ALUCtrl.scala 94:31]
  wire  _T_41 = 32'h1003 == _T; // @[ALUCtrl.scala 95:31]
  wire  _T_43 = 32'h2003 == _T; // @[ALUCtrl.scala 96:31]
  wire  _T_47 = 32'h5003 == _T; // @[ALUCtrl.scala 98:31]
  wire  _T_49 = 32'h6003 == _T; // @[ALUCtrl.scala 99:31]
  wire  _T_51 = 32'h3 == _T; // @[ALUCtrl.scala 100:31]
  wire  _T_53 = 32'h6013 == _T; // @[ALUCtrl.scala 101:31]
  wire  _T_55 = 32'h3033 == _T_22; // @[ALUCtrl.scala 102:31]
  wire  _T_57 = 32'h3b == _T_22; // @[ALUCtrl.scala 103:31]
  wire  _T_59 = 32'h4000003b == _T_22; // @[ALUCtrl.scala 104:31]
  wire  _T_61 = 32'h7033 == _T_22; // @[ALUCtrl.scala 105:31]
  wire  _T_63 = 32'h33 == _T_22; // @[ALUCtrl.scala 106:31]
  wire  _T_65 = 32'h200503b == _T_22; // @[ALUCtrl.scala 107:31]
  wire  _T_67 = 32'h200703b == _T_22; // @[ALUCtrl.scala 108:31]
  wire  _T_69 = 32'h40000033 == _T_22; // @[ALUCtrl.scala 109:31]
  wire  _T_71 = 32'h200003b == _T_22; // @[ALUCtrl.scala 110:31]
  wire  _T_73 = 32'h200603b == _T_22; // @[ALUCtrl.scala 111:31]
  wire  _T_75 = 32'h200403b == _T_22; // @[ALUCtrl.scala 112:31]
  wire  _T_77 = 32'h2000033 == _T_22; // @[ALUCtrl.scala 113:31]
  wire  _T_79 = 32'h6033 == _T_22; // @[ALUCtrl.scala 114:31]
  wire  _T_81 = 32'h103b == _T_22; // @[ALUCtrl.scala 115:31]
  wire  _T_83 = 32'h4000503b == _T_22; // @[ALUCtrl.scala 116:31]
  wire  _T_85 = 32'h503b == _T_22; // @[ALUCtrl.scala 117:31]
  wire  _T_87 = 32'h2033 == _T_22; // @[ALUCtrl.scala 118:31]
  wire  _T_89 = 32'h2005033 == _T_22; // @[ALUCtrl.scala 119:31]
  wire  _T_91 = 32'h4033 == _T_22; // @[ALUCtrl.scala 120:31]
  wire  _T_93 = 32'h2006033 == _T_22; // @[ALUCtrl.scala 121:31]
  wire  _T_95 = 32'h2004033 == _T_22; // @[ALUCtrl.scala 122:31]
  wire  _T_97 = 32'h1033 == _T_22; // @[ALUCtrl.scala 123:31]
  wire  _T_99 = 32'h63 == _T; // @[ALUCtrl.scala 124:31]
  wire  _T_101 = 32'h6063 == _T; // @[ALUCtrl.scala 125:31]
  wire  _T_103 = 32'h7063 == _T; // @[ALUCtrl.scala 126:31]
  wire  _T_105 = 32'h4063 == _T; // @[ALUCtrl.scala 127:31]
  wire  _T_107 = 32'h5063 == _T; // @[ALUCtrl.scala 128:31]
  wire  _T_109 = 32'h1063 == _T; // @[ALUCtrl.scala 129:31]
  wire  _T_111 = 32'h2007033 == _T_22; // @[ALUCtrl.scala 130:31]
  wire  _T_113 = 32'h5033 == _T_22; // @[ALUCtrl.scala 131:31]
  wire [4:0] _io_ALUCtrl_T = _T_113 ? 5'h8 : 5'h1f; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_1 = _T_111 ? 5'h1d : _io_ALUCtrl_T; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_2 = _T_109 ? 5'hb : _io_ALUCtrl_T_1; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_3 = _T_107 ? 5'h1c : _io_ALUCtrl_T_2; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_4 = _T_105 ? 5'h5 : _io_ALUCtrl_T_3; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_5 = _T_103 ? 5'h1b : _io_ALUCtrl_T_4; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_6 = _T_101 ? 5'h7 : _io_ALUCtrl_T_5; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_7 = _T_99 ? 5'h1a : _io_ALUCtrl_T_6; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_8 = _T_97 ? 5'h6 : _io_ALUCtrl_T_7; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_9 = _T_95 ? 5'h19 : _io_ALUCtrl_T_8; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_10 = _T_93 ? 5'h18 : _io_ALUCtrl_T_9; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_11 = _T_91 ? 5'h4 : _io_ALUCtrl_T_10; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_12 = _T_89 ? 5'h17 : _io_ALUCtrl_T_11; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_13 = _T_87 ? 5'h5 : _io_ALUCtrl_T_12; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_14 = _T_85 ? 5'hc : _io_ALUCtrl_T_13; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_15 = _T_83 ? 5'hf : _io_ALUCtrl_T_14; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_16 = _T_81 ? 5'he : _io_ALUCtrl_T_15; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_17 = _T_79 ? 5'h3 : _io_ALUCtrl_T_16; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_18 = _T_77 ? 5'h16 : _io_ALUCtrl_T_17; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_19 = _T_75 ? 5'h15 : _io_ALUCtrl_T_18; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_20 = _T_73 ? 5'h14 : _io_ALUCtrl_T_19; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_21 = _T_71 ? 5'h13 : _io_ALUCtrl_T_20; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_22 = _T_69 ? 5'h1 : _io_ALUCtrl_T_21; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_23 = _T_67 ? 5'h12 : _io_ALUCtrl_T_22; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_24 = _T_65 ? 5'h11 : _io_ALUCtrl_T_23; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_25 = _T_63 ? 5'h0 : _io_ALUCtrl_T_24; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_26 = _T_61 ? 5'h2 : _io_ALUCtrl_T_25; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_27 = _T_59 ? 5'h10 : _io_ALUCtrl_T_26; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_28 = _T_57 ? 5'hd : _io_ALUCtrl_T_27; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_29 = _T_55 ? 5'h7 : _io_ALUCtrl_T_28; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_30 = _T_53 ? 5'h3 : _io_ALUCtrl_T_29; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_31 = _T_51 ? 5'h0 : _io_ALUCtrl_T_30; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_32 = _T_49 ? 5'h0 : _io_ALUCtrl_T_31; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_33 = _T_47 ? 5'h0 : _io_ALUCtrl_T_32; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_34 = _T_17 ? 5'h0 : _io_ALUCtrl_T_33; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_35 = _T_43 ? 5'h0 : _io_ALUCtrl_T_34; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_36 = _T_41 ? 5'h0 : _io_ALUCtrl_T_35; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_37 = _T_39 ? 5'h9 : _io_ALUCtrl_T_36; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_38 = _T_37 ? 5'hf : _io_ALUCtrl_T_37; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_39 = _T_35 ? 5'he : _io_ALUCtrl_T_38; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_40 = _T_33 ? 5'h8 : _io_ALUCtrl_T_39; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_41 = _T_31 ? 5'hd : _io_ALUCtrl_T_40; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_42 = _T_29 ? 5'h4 : _io_ALUCtrl_T_41; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_43 = _T_27 ? 5'h2 : _io_ALUCtrl_T_42; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_44 = _T_25 ? 5'h6 : _io_ALUCtrl_T_43; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_45 = _T_23 ? 5'hc : _io_ALUCtrl_T_44; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_46 = _T_21 ? 5'h7 : _io_ALUCtrl_T_45; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_47 = _T_19 ? 5'h0 : _io_ALUCtrl_T_46; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_48 = _T_17 ? 5'h0 : _io_ALUCtrl_T_47; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_49 = _T_15 ? 5'h1f : _io_ALUCtrl_T_48; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_50 = _T_13 ? 5'h0 : _io_ALUCtrl_T_49; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_51 = _T_11 ? 5'ha : _io_ALUCtrl_T_50; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_52 = _T_9 ? 5'h0 : _io_ALUCtrl_T_51; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_53 = _T_7 ? 5'h0 : _io_ALUCtrl_T_52; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_54 = _T_5 ? 5'h0 : _io_ALUCtrl_T_53; // @[Mux.scala 98:16]
  wire [4:0] _io_ALUCtrl_T_55 = _T_3 ? 5'h0 : _io_ALUCtrl_T_54; // @[Mux.scala 98:16]
  assign io_ALUCtrl = _T_1 ? 5'h0 : _io_ALUCtrl_T_55; // @[Mux.scala 98:16]
endmodule
module ALUSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_AluSrc1,
  output [1:0]  io_AluSrc2
);
  wire [31:0] _T = io_inst & 32'hfc00707f; // @[ALUSrcGen.scala 63:49]
  wire  _T_1 = 32'h1013 == _T; // @[ALUSrcGen.scala 63:49]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[ALUSrcGen.scala 63:49]
  wire  _T_3 = 32'h13 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire [31:0] _T_4 = io_inst & 32'hfe00707f; // @[ALUSrcGen.scala 63:49]
  wire  _T_5 = 32'h101b == _T_4; // @[ALUSrcGen.scala 63:49]
  wire  _T_7 = 32'h5013 == _T; // @[ALUSrcGen.scala 63:49]
  wire  _T_9 = 32'h6063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_11 = 32'h6013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_13 = 32'h7013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_15 = 32'h4063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_17 = 32'h2007033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_19 = 32'h503b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_21 = 32'h501b == _T_4; // @[ALUSrcGen.scala 63:49]
  wire  _T_23 = 32'h3003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_25 = 32'h3013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_27 = 32'h3b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_29 = 32'h2000033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_31 = 32'h7033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_33 = 32'h103b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_35 = 32'h1003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_37 = 32'h200603b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_39 = 32'h3033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_41 = 32'h2033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_43 = 32'h200403b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_45 = 32'h4000501b == _T_4; // @[ALUSrcGen.scala 63:49]
  wire  _T_47 = 32'h1033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_49 = 32'h67 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_51 = 32'h4000503b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_53 = 32'h1063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_55 = 32'h1b == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_57 = 32'h3023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_59 = 32'h200503b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_61 = 32'h4013 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_63 = 32'h2003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_65 = 32'h4003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_67 = 32'h2005033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_69 = 32'h4000003b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_71 = 32'h5003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_73 = 32'h3 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_75 = 32'h7063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_77 = 32'h23 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_79 = 32'h33 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_81 = 32'h2023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire  _T_83 = 32'h6033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_85 = 32'h2004033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_87 = 32'h4033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_89 = 32'h40005013 == _T; // @[ALUSrcGen.scala 63:49]
  wire  _T_91 = 32'h63 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_93 = 32'h40000033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_95 = 32'h5033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_97 = 32'h5063 == _T_2; // @[ALUSrcGen.scala 65:49]
  wire  _T_99 = 32'h200703b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_101 = 32'h6003 == _T_2; // @[ALUSrcGen.scala 63:49]
  wire  _T_103 = 32'h200003b == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_105 = 32'h2006033 == _T_4; // @[ALUSrcGen.scala 66:49]
  wire  _T_107 = 32'h1023 == _T_2; // @[ALUSrcGen.scala 64:49]
  wire [31:0] _T_108 = io_inst & 32'h7f; // @[ALUSrcGen.scala 71:31]
  wire  _T_109 = 32'h17 == _T_108; // @[ALUSrcGen.scala 71:31]
  wire  _T_111 = 32'h37 == _T_108; // @[ALUSrcGen.scala 72:31]
  wire  _io_AluSrc1_T_2 = _T_107 ? 1'h0 : _T_109 | _T_111; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_3 = _T_105 ? 1'h0 : _io_AluSrc1_T_2; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_4 = _T_103 ? 1'h0 : _io_AluSrc1_T_3; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_5 = _T_101 ? 1'h0 : _io_AluSrc1_T_4; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_6 = _T_99 ? 1'h0 : _io_AluSrc1_T_5; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_7 = _T_97 ? 1'h0 : _io_AluSrc1_T_6; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_8 = _T_95 ? 1'h0 : _io_AluSrc1_T_7; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_9 = _T_93 ? 1'h0 : _io_AluSrc1_T_8; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_10 = _T_91 ? 1'h0 : _io_AluSrc1_T_9; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_11 = _T_89 ? 1'h0 : _io_AluSrc1_T_10; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_12 = _T_87 ? 1'h0 : _io_AluSrc1_T_11; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_13 = _T_85 ? 1'h0 : _io_AluSrc1_T_12; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_14 = _T_83 ? 1'h0 : _io_AluSrc1_T_13; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_15 = _T_81 ? 1'h0 : _io_AluSrc1_T_14; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_16 = _T_79 ? 1'h0 : _io_AluSrc1_T_15; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_17 = _T_77 ? 1'h0 : _io_AluSrc1_T_16; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_18 = _T_75 ? 1'h0 : _io_AluSrc1_T_17; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_19 = _T_73 ? 1'h0 : _io_AluSrc1_T_18; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_20 = _T_71 ? 1'h0 : _io_AluSrc1_T_19; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_21 = _T_69 ? 1'h0 : _io_AluSrc1_T_20; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_22 = _T_67 ? 1'h0 : _io_AluSrc1_T_21; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_23 = _T_65 ? 1'h0 : _io_AluSrc1_T_22; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_24 = _T_63 ? 1'h0 : _io_AluSrc1_T_23; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_25 = _T_61 ? 1'h0 : _io_AluSrc1_T_24; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_26 = _T_59 ? 1'h0 : _io_AluSrc1_T_25; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_27 = _T_57 ? 1'h0 : _io_AluSrc1_T_26; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_28 = _T_55 ? 1'h0 : _io_AluSrc1_T_27; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_29 = _T_53 ? 1'h0 : _io_AluSrc1_T_28; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_30 = _T_51 ? 1'h0 : _io_AluSrc1_T_29; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_31 = _T_49 ? 1'h0 : _io_AluSrc1_T_30; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_32 = _T_47 ? 1'h0 : _io_AluSrc1_T_31; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_33 = _T_45 ? 1'h0 : _io_AluSrc1_T_32; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_34 = _T_43 ? 1'h0 : _io_AluSrc1_T_33; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_35 = _T_41 ? 1'h0 : _io_AluSrc1_T_34; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_36 = _T_39 ? 1'h0 : _io_AluSrc1_T_35; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_37 = _T_37 ? 1'h0 : _io_AluSrc1_T_36; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_38 = _T_35 ? 1'h0 : _io_AluSrc1_T_37; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_39 = _T_33 ? 1'h0 : _io_AluSrc1_T_38; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_40 = _T_31 ? 1'h0 : _io_AluSrc1_T_39; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_41 = _T_29 ? 1'h0 : _io_AluSrc1_T_40; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_42 = _T_27 ? 1'h0 : _io_AluSrc1_T_41; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_43 = _T_25 ? 1'h0 : _io_AluSrc1_T_42; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_44 = _T_23 ? 1'h0 : _io_AluSrc1_T_43; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_45 = _T_21 ? 1'h0 : _io_AluSrc1_T_44; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_46 = _T_19 ? 1'h0 : _io_AluSrc1_T_45; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_47 = _T_17 ? 1'h0 : _io_AluSrc1_T_46; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_48 = _T_15 ? 1'h0 : _io_AluSrc1_T_47; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_49 = _T_13 ? 1'h0 : _io_AluSrc1_T_48; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_50 = _T_11 ? 1'h0 : _io_AluSrc1_T_49; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_51 = _T_9 ? 1'h0 : _io_AluSrc1_T_50; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_52 = _T_7 ? 1'h0 : _io_AluSrc1_T_51; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_53 = _T_5 ? 1'h0 : _io_AluSrc1_T_52; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_54 = _T_3 ? 1'h0 : _io_AluSrc1_T_53; // @[Mux.scala 98:16]
  wire  _io_AluSrc1_T_55 = _T_1 ? 1'h0 : _io_AluSrc1_T_54; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T = _T_111 ? 2'h3 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_1 = _T_109 ? 2'h2 : _io_AluSrc2_T; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_2 = _T_107 ? 2'h1 : _io_AluSrc2_T_1; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_3 = _T_105 ? 2'h0 : _io_AluSrc2_T_2; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_4 = _T_103 ? 2'h0 : _io_AluSrc2_T_3; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_5 = _T_101 ? 2'h1 : _io_AluSrc2_T_4; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_6 = _T_99 ? 2'h0 : _io_AluSrc2_T_5; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_7 = _T_97 ? 2'h0 : _io_AluSrc2_T_6; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_8 = _T_95 ? 2'h0 : _io_AluSrc2_T_7; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_9 = _T_93 ? 2'h0 : _io_AluSrc2_T_8; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_10 = _T_91 ? 2'h0 : _io_AluSrc2_T_9; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_11 = _T_89 ? 2'h1 : _io_AluSrc2_T_10; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_12 = _T_87 ? 2'h0 : _io_AluSrc2_T_11; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_13 = _T_85 ? 2'h0 : _io_AluSrc2_T_12; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_14 = _T_83 ? 2'h0 : _io_AluSrc2_T_13; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_15 = _T_81 ? 2'h1 : _io_AluSrc2_T_14; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_16 = _T_79 ? 2'h0 : _io_AluSrc2_T_15; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_17 = _T_77 ? 2'h1 : _io_AluSrc2_T_16; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_18 = _T_75 ? 2'h0 : _io_AluSrc2_T_17; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_19 = _T_73 ? 2'h1 : _io_AluSrc2_T_18; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_20 = _T_71 ? 2'h1 : _io_AluSrc2_T_19; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_21 = _T_69 ? 2'h0 : _io_AluSrc2_T_20; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_22 = _T_67 ? 2'h0 : _io_AluSrc2_T_21; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_23 = _T_65 ? 2'h1 : _io_AluSrc2_T_22; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_24 = _T_63 ? 2'h1 : _io_AluSrc2_T_23; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_25 = _T_61 ? 2'h1 : _io_AluSrc2_T_24; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_26 = _T_59 ? 2'h0 : _io_AluSrc2_T_25; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_27 = _T_57 ? 2'h1 : _io_AluSrc2_T_26; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_28 = _T_55 ? 2'h1 : _io_AluSrc2_T_27; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_29 = _T_53 ? 2'h0 : _io_AluSrc2_T_28; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_30 = _T_51 ? 2'h0 : _io_AluSrc2_T_29; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_31 = _T_49 ? 2'h1 : _io_AluSrc2_T_30; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_32 = _T_47 ? 2'h0 : _io_AluSrc2_T_31; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_33 = _T_45 ? 2'h1 : _io_AluSrc2_T_32; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_34 = _T_43 ? 2'h0 : _io_AluSrc2_T_33; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_35 = _T_41 ? 2'h0 : _io_AluSrc2_T_34; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_36 = _T_39 ? 2'h0 : _io_AluSrc2_T_35; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_37 = _T_37 ? 2'h0 : _io_AluSrc2_T_36; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_38 = _T_35 ? 2'h1 : _io_AluSrc2_T_37; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_39 = _T_33 ? 2'h0 : _io_AluSrc2_T_38; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_40 = _T_31 ? 2'h0 : _io_AluSrc2_T_39; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_41 = _T_29 ? 2'h0 : _io_AluSrc2_T_40; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_42 = _T_27 ? 2'h0 : _io_AluSrc2_T_41; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_43 = _T_25 ? 2'h1 : _io_AluSrc2_T_42; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_44 = _T_23 ? 2'h1 : _io_AluSrc2_T_43; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_45 = _T_21 ? 2'h1 : _io_AluSrc2_T_44; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_46 = _T_19 ? 2'h0 : _io_AluSrc2_T_45; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_47 = _T_17 ? 2'h0 : _io_AluSrc2_T_46; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_48 = _T_15 ? 2'h0 : _io_AluSrc2_T_47; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_49 = _T_13 ? 2'h1 : _io_AluSrc2_T_48; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_50 = _T_11 ? 2'h1 : _io_AluSrc2_T_49; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_51 = _T_9 ? 2'h0 : _io_AluSrc2_T_50; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_52 = _T_7 ? 2'h1 : _io_AluSrc2_T_51; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_53 = _T_5 ? 2'h1 : _io_AluSrc2_T_52; // @[Mux.scala 98:16]
  wire [1:0] _io_AluSrc2_T_54 = _T_3 ? 2'h1 : _io_AluSrc2_T_53; // @[Mux.scala 98:16]
  assign io_AluSrc1 = {{1'd0}, _io_AluSrc1_T_55}; // @[Mux.scala 98:16]
  assign io_AluSrc2 = _T_1 ? 2'h1 : _io_AluSrc2_T_54; // @[Mux.scala 98:16]
endmodule
module memWriteMGen(
  input  [31:0] io_inst,
  output        io_memWriteM
);
  wire [31:0] _T = io_inst & 32'h707f; // @[memWriteMGen.scala 19:49]
  wire  _T_1 = 32'h3023 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_3 = 32'h23 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_5 = 32'h2023 == _T; // @[memWriteMGen.scala 19:49]
  wire  _T_7 = 32'h1023 == _T; // @[memWriteMGen.scala 19:49]
  assign io_memWriteM = _T_1 | (_T_3 | (_T_5 | _T_7)); // @[Mux.scala 98:16]
endmodule
module memWriteMaskGen(
  input  [31:0] io_inst,
  output [7:0]  io_mask
);
  wire [7:0] _io_mask_T_2 = 3'h0 == io_inst[14:12] ? 8'h1 : 8'h0; // @[Mux.scala 80:57]
  wire [7:0] _io_mask_T_4 = 3'h1 == io_inst[14:12] ? 8'h3 : _io_mask_T_2; // @[Mux.scala 80:57]
  wire [7:0] _io_mask_T_6 = 3'h2 == io_inst[14:12] ? 8'hf : _io_mask_T_4; // @[Mux.scala 80:57]
  assign io_mask = 3'h3 == io_inst[14:12] ? 8'hff : _io_mask_T_6; // @[Mux.scala 80:57]
endmodule
module memReadNumGen(
  input  [31:0] io_inst,
  output [2:0]  io_memReadNum
);
  assign io_memReadNum = io_inst[14:12]; // @[instDe.scala 13:16]
endmodule
module dnpcSrcGen(
  input  [31:0] io_inst,
  output        io_dnpcSrc
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 25:49]
  wire  _T_1 = 32'h6063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_3 = 32'h4063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_5 = 32'h1063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_7 = 32'h7063 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_9 = 32'h63 == _T; // @[npcSrcGen.scala 25:49]
  wire  _T_11 = 32'h5063 == _T; // @[npcSrcGen.scala 25:49]
  wire [31:0] _T_12 = io_inst & 32'h7f; // @[npcSrcGen.scala 30:31]
  wire  _T_13 = 32'h6f == _T_12; // @[npcSrcGen.scala 30:31]
  assign io_dnpcSrc = _T_1 | (_T_3 | (_T_5 | (_T_7 | (_T_9 | (_T_11 | _T_13))))); // @[Mux.scala 98:16]
endmodule
module jumpGen(
  input  [31:0] io_inst,
  output        io_jump
);
  wire [31:0] _T = io_inst & 32'h7f; // @[npcSrcGen.scala 46:14]
  wire  _T_1 = 32'h6f == _T; // @[npcSrcGen.scala 46:14]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[npcSrcGen.scala 47:14]
  wire  _T_3 = 32'h67 == _T_2; // @[npcSrcGen.scala 47:14]
  assign io_jump = _T_1 | _T_3; // @[Mux.scala 98:16]
endmodule
module branchGen(
  input  [31:0] io_inst,
  output        io_branch
);
  wire [31:0] _T = io_inst & 32'h707f; // @[npcSrcGen.scala 66:47]
  wire  _T_1 = 32'h6063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_3 = 32'h4063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_5 = 32'h1063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_7 = 32'h7063 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_9 = 32'h63 == _T; // @[npcSrcGen.scala 66:47]
  wire  _T_11 = 32'h5063 == _T; // @[npcSrcGen.scala 66:47]
  assign io_branch = _T_1 | (_T_3 | (_T_5 | (_T_7 | (_T_9 | _T_11)))); // @[Mux.scala 98:16]
endmodule
module regEnGen(
  input  [31:0] io_inst,
  output        io_regEn
);
  wire [31:0] _T = io_inst & 32'hfc00707f; // @[regEnGen.scala 33:45]
  wire  _T_1 = 32'h1013 == _T; // @[regEnGen.scala 33:45]
  wire [31:0] _T_2 = io_inst & 32'h707f; // @[regEnGen.scala 33:45]
  wire  _T_3 = 32'h13 == _T_2; // @[regEnGen.scala 33:45]
  wire [31:0] _T_4 = io_inst & 32'hfe00707f; // @[regEnGen.scala 33:45]
  wire  _T_5 = 32'h101b == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_7 = 32'h5013 == _T; // @[regEnGen.scala 33:45]
  wire  _T_9 = 32'h6063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_11 = 32'h6013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_13 = 32'h7013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_15 = 32'h4063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_17 = 32'h2007033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_19 = 32'h503b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_21 = 32'h501b == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_23 = 32'h3003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_25 = 32'h3013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_27 = 32'h3b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_29 = 32'h2000033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_31 = 32'h7033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_33 = 32'h103b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_35 = 32'h1003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_37 = 32'h200603b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_39 = 32'h3033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_41 = 32'h2033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_43 = 32'h200403b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_45 = 32'h4000501b == _T_4; // @[regEnGen.scala 33:45]
  wire  _T_47 = 32'h1033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_49 = 32'h67 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_51 = 32'h4000503b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_53 = 32'h1063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_55 = 32'h1b == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_57 = 32'h3023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_59 = 32'h200503b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_61 = 32'h4013 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_63 = 32'h2003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_65 = 32'h4003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_67 = 32'h2005033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_69 = 32'h4000003b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_71 = 32'h5003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_73 = 32'h3 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_75 = 32'h7063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_77 = 32'h23 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_79 = 32'h33 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_81 = 32'h2023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_83 = 32'h6033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_85 = 32'h2004033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_87 = 32'h4033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_89 = 32'h40005013 == _T; // @[regEnGen.scala 33:45]
  wire  _T_91 = 32'h63 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_93 = 32'h40000033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_95 = 32'h5033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_97 = 32'h5063 == _T_2; // @[regEnGen.scala 37:45]
  wire  _T_99 = 32'h200703b == _T_4; // @[regEnGen.scala 35:45]
  wire [31:0] _T_100 = io_inst & 32'h7f; // @[regEnGen.scala 32:45]
  wire  _T_101 = 32'h17 == _T_100; // @[regEnGen.scala 32:45]
  wire  _T_103 = 32'h6003 == _T_2; // @[regEnGen.scala 33:45]
  wire  _T_105 = 32'h200003b == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_107 = 32'h37 == _T_100; // @[regEnGen.scala 32:45]
  wire  _T_109 = 32'h2006033 == _T_4; // @[regEnGen.scala 35:45]
  wire  _T_111 = 32'h1023 == _T_2; // @[regEnGen.scala 36:45]
  wire  _T_113 = 32'h6f == _T_100; // @[regEnGen.scala 34:45]
  wire  _io_regEn_T_1 = _T_111 ? 1'h0 : _T_113; // @[Mux.scala 98:16]
  wire  _io_regEn_T_8 = _T_97 ? 1'h0 : _T_99 | (_T_101 | (_T_103 | (_T_105 | (_T_107 | (_T_109 | _io_regEn_T_1))))); // @[Mux.scala 98:16]
  wire  _io_regEn_T_11 = _T_91 ? 1'h0 : _T_93 | (_T_95 | _io_regEn_T_8); // @[Mux.scala 98:16]
  wire  _io_regEn_T_16 = _T_81 ? 1'h0 : _T_83 | (_T_85 | (_T_87 | (_T_89 | _io_regEn_T_11))); // @[Mux.scala 98:16]
  wire  _io_regEn_T_18 = _T_77 ? 1'h0 : _T_79 | _io_regEn_T_16; // @[Mux.scala 98:16]
  wire  _io_regEn_T_19 = _T_75 ? 1'h0 : _io_regEn_T_18; // @[Mux.scala 98:16]
  wire  _io_regEn_T_28 = _T_57 ? 1'h0 : _T_59 | (_T_61 | (_T_63 | (_T_65 | (_T_67 | (_T_69 | (_T_71 | (_T_73 |
    _io_regEn_T_19))))))); // @[Mux.scala 98:16]
  wire  _io_regEn_T_30 = _T_53 ? 1'h0 : _T_55 | _io_regEn_T_28; // @[Mux.scala 98:16]
  wire  _io_regEn_T_49 = _T_15 ? 1'h0 : _T_17 | (_T_19 | (_T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29 | (_T_31 | (_T_33 |
    (_T_35 | (_T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | _io_regEn_T_30))))))))))))))))); // @[Mux.scala 98:16]
  wire  _io_regEn_T_52 = _T_9 ? 1'h0 : _T_11 | (_T_13 | _io_regEn_T_49); // @[Mux.scala 98:16]
  assign io_regEn = _T_1 | (_T_3 | (_T_5 | (_T_7 | _io_regEn_T_52))); // @[Mux.scala 98:16]
endmodule
module ResultSrcGen(
  input  [31:0] io_inst,
  output [1:0]  io_ResultSrc
);
  wire [31:0] _T = io_inst & 32'hfe00707f; // @[ResultSrcGen.scala 39:44]
  wire  _T_1 = 32'h2007033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_3 = 32'h503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_5 = 32'h3b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_7 = 32'h2000033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_9 = 32'h7033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_11 = 32'h103b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_13 = 32'h200603b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_15 = 32'h3033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_17 = 32'h2033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_19 = 32'h200403b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_21 = 32'h1033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_23 = 32'h4000503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_25 = 32'h200503b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_27 = 32'h2005033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_29 = 32'h4000003b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_31 = 32'h33 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_33 = 32'h6033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_35 = 32'h2004033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_37 = 32'h4033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_39 = 32'h40000033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_41 = 32'h5033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_43 = 32'h200703b == _T; // @[ResultSrcGen.scala 39:44]
  wire [31:0] _T_44 = io_inst & 32'h7f; // @[ResultSrcGen.scala 37:44]
  wire  _T_45 = 32'h17 == _T_44; // @[ResultSrcGen.scala 37:44]
  wire  _T_47 = 32'h200003b == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_49 = 32'h37 == _T_44; // @[ResultSrcGen.scala 37:44]
  wire  _T_51 = 32'h2006033 == _T; // @[ResultSrcGen.scala 39:44]
  wire  _T_53 = 32'h6f == _T_44; // @[ResultSrcGen.scala 38:44]
  wire [31:0] _T_54 = io_inst & 32'h707f; // @[ResultSrcGen.scala 44:26]
  wire  _T_55 = 32'h13 == _T_54; // @[ResultSrcGen.scala 44:26]
  wire  _T_57 = 32'h67 == _T_54; // @[ResultSrcGen.scala 45:26]
  wire  _T_61 = 32'h3003 == _T_54; // @[ResultSrcGen.scala 47:26]
  wire  _T_63 = 32'h4003 == _T_54; // @[ResultSrcGen.scala 48:26]
  wire  _T_65 = 32'h3013 == _T_54; // @[ResultSrcGen.scala 49:26]
  wire  _T_67 = 32'h501b == _T; // @[ResultSrcGen.scala 50:26]
  wire [31:0] _T_68 = io_inst & 32'hfc00707f; // @[ResultSrcGen.scala 51:26]
  wire  _T_69 = 32'h1013 == _T_68; // @[ResultSrcGen.scala 51:26]
  wire  _T_71 = 32'h7013 == _T_54; // @[ResultSrcGen.scala 52:26]
  wire  _T_73 = 32'h4013 == _T_54; // @[ResultSrcGen.scala 53:26]
  wire  _T_75 = 32'h1b == _T_54; // @[ResultSrcGen.scala 54:26]
  wire  _T_77 = 32'h5013 == _T_68; // @[ResultSrcGen.scala 55:26]
  wire  _T_79 = 32'h101b == _T; // @[ResultSrcGen.scala 56:26]
  wire  _T_81 = 32'h4000501b == _T; // @[ResultSrcGen.scala 57:26]
  wire  _T_83 = 32'h40005013 == _T_68; // @[ResultSrcGen.scala 58:26]
  wire  _T_85 = 32'h6013 == _T_54; // @[ResultSrcGen.scala 59:26]
  wire  _T_87 = 32'h1003 == _T_54; // @[ResultSrcGen.scala 60:26]
  wire  _T_89 = 32'h2003 == _T_54; // @[ResultSrcGen.scala 61:26]
  wire  _T_91 = 32'h5003 == _T_54; // @[ResultSrcGen.scala 62:26]
  wire  _T_93 = 32'h6003 == _T_54; // @[ResultSrcGen.scala 63:26]
  wire  _T_95 = 32'h3 == _T_54; // @[ResultSrcGen.scala 64:26]
  wire [1:0] _io_ResultSrc_T_2 = _T_95 ? 2'h2 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_3 = _T_93 ? 2'h2 : _io_ResultSrc_T_2; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_4 = _T_91 ? 2'h2 : _io_ResultSrc_T_3; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_5 = _T_89 ? 2'h2 : _io_ResultSrc_T_4; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_6 = _T_87 ? 2'h2 : _io_ResultSrc_T_5; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_7 = _T_85 ? 2'h0 : _io_ResultSrc_T_6; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_8 = _T_83 ? 2'h0 : _io_ResultSrc_T_7; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_9 = _T_81 ? 2'h0 : _io_ResultSrc_T_8; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_10 = _T_79 ? 2'h0 : _io_ResultSrc_T_9; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_11 = _T_77 ? 2'h0 : _io_ResultSrc_T_10; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_12 = _T_75 ? 2'h0 : _io_ResultSrc_T_11; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_13 = _T_73 ? 2'h0 : _io_ResultSrc_T_12; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_14 = _T_71 ? 2'h0 : _io_ResultSrc_T_13; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_15 = _T_69 ? 2'h0 : _io_ResultSrc_T_14; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_16 = _T_67 ? 2'h0 : _io_ResultSrc_T_15; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_17 = _T_65 ? 2'h0 : _io_ResultSrc_T_16; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_18 = _T_63 ? 2'h2 : _io_ResultSrc_T_17; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_19 = _T_61 ? 2'h2 : _io_ResultSrc_T_18; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_20 = _T_57 ? 2'h1 : _io_ResultSrc_T_19; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_21 = _T_57 ? 2'h1 : _io_ResultSrc_T_20; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_22 = _T_55 ? 2'h0 : _io_ResultSrc_T_21; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_23 = _T_53 ? 2'h1 : _io_ResultSrc_T_22; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_24 = _T_51 ? 2'h0 : _io_ResultSrc_T_23; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_25 = _T_49 ? 2'h0 : _io_ResultSrc_T_24; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_26 = _T_47 ? 2'h0 : _io_ResultSrc_T_25; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_27 = _T_45 ? 2'h0 : _io_ResultSrc_T_26; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_28 = _T_43 ? 2'h0 : _io_ResultSrc_T_27; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_29 = _T_41 ? 2'h0 : _io_ResultSrc_T_28; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_30 = _T_39 ? 2'h0 : _io_ResultSrc_T_29; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_31 = _T_37 ? 2'h0 : _io_ResultSrc_T_30; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_32 = _T_35 ? 2'h0 : _io_ResultSrc_T_31; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_33 = _T_33 ? 2'h0 : _io_ResultSrc_T_32; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_34 = _T_31 ? 2'h0 : _io_ResultSrc_T_33; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_35 = _T_29 ? 2'h0 : _io_ResultSrc_T_34; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_36 = _T_27 ? 2'h0 : _io_ResultSrc_T_35; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_37 = _T_25 ? 2'h0 : _io_ResultSrc_T_36; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_38 = _T_23 ? 2'h0 : _io_ResultSrc_T_37; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_39 = _T_21 ? 2'h0 : _io_ResultSrc_T_38; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_40 = _T_19 ? 2'h0 : _io_ResultSrc_T_39; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_41 = _T_17 ? 2'h0 : _io_ResultSrc_T_40; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_42 = _T_15 ? 2'h0 : _io_ResultSrc_T_41; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_43 = _T_13 ? 2'h0 : _io_ResultSrc_T_42; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_44 = _T_11 ? 2'h0 : _io_ResultSrc_T_43; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_45 = _T_9 ? 2'h0 : _io_ResultSrc_T_44; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_46 = _T_7 ? 2'h0 : _io_ResultSrc_T_45; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_47 = _T_5 ? 2'h0 : _io_ResultSrc_T_46; // @[Mux.scala 98:16]
  wire [1:0] _io_ResultSrc_T_48 = _T_3 ? 2'h0 : _io_ResultSrc_T_47; // @[Mux.scala 98:16]
  assign io_ResultSrc = _T_1 ? 2'h0 : _io_ResultSrc_T_48; // @[Mux.scala 98:16]
endmodule
module CtrlUnit(
  input  [31:0] io_inst,
  output [1:0]  io_CtrlS_AluSrc1,
  output [1:0]  io_CtrlS_AluSrc2,
  output [4:0]  io_CtrlS_ALUCtrl,
  output        io_CtrlS_memWriteM,
  output [7:0]  io_CtrlS_memWriteMask,
  output [2:0]  io_CtrlS_memReadNum,
  output        io_CtrlS_dnpcSrc,
  output        io_CtrlS_jump,
  output        io_CtrlS_branch,
  output        io_CtrlS_regEn,
  output [1:0]  io_CtrlS_ResultSrc,
  output        io_CtrlS_fencei
);
  wire [31:0] ALUCtrl_ins_io_inst; // @[CtrlUnit.scala 33:26]
  wire [4:0] ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 33:26]
  wire [31:0] ALUSrcGen_ins_io_inst; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 37:29]
  wire [1:0] ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 37:29]
  wire [31:0] memWriteMGen_ins_io_inst; // @[CtrlUnit.scala 42:32]
  wire  memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 42:32]
  wire [31:0] memWriteMaskGen_ins_io_inst; // @[CtrlUnit.scala 46:35]
  wire [7:0] memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 46:35]
  wire [31:0] memReadNumGen_ins_io_inst; // @[CtrlUnit.scala 50:33]
  wire [2:0] memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 50:33]
  wire [31:0] dnpcSrcGen_ins_io_inst; // @[CtrlUnit.scala 54:32]
  wire  dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 54:32]
  wire [31:0] jumpGen_ins_io_inst; // @[CtrlUnit.scala 58:27]
  wire  jumpGen_ins_io_jump; // @[CtrlUnit.scala 58:27]
  wire [31:0] branchGen_ins_io_inst; // @[CtrlUnit.scala 62:29]
  wire  branchGen_ins_io_branch; // @[CtrlUnit.scala 62:29]
  wire [31:0] regEnGen_ins_io_inst; // @[CtrlUnit.scala 67:28]
  wire  regEnGen_ins_io_regEn; // @[CtrlUnit.scala 67:28]
  wire [31:0] ResultSrcGen_ins_io_inst; // @[CtrlUnit.scala 71:32]
  wire [1:0] ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 71:32]
  wire [31:0] _io_CtrlS_fencei_T = io_inst & 32'h707f; // @[CtrlUnit.scala 75:30]
  ALUCtrl ALUCtrl_ins ( // @[CtrlUnit.scala 33:26]
    .io_inst(ALUCtrl_ins_io_inst),
    .io_ALUCtrl(ALUCtrl_ins_io_ALUCtrl)
  );
  ALUSrcGen ALUSrcGen_ins ( // @[CtrlUnit.scala 37:29]
    .io_inst(ALUSrcGen_ins_io_inst),
    .io_AluSrc1(ALUSrcGen_ins_io_AluSrc1),
    .io_AluSrc2(ALUSrcGen_ins_io_AluSrc2)
  );
  memWriteMGen memWriteMGen_ins ( // @[CtrlUnit.scala 42:32]
    .io_inst(memWriteMGen_ins_io_inst),
    .io_memWriteM(memWriteMGen_ins_io_memWriteM)
  );
  memWriteMaskGen memWriteMaskGen_ins ( // @[CtrlUnit.scala 46:35]
    .io_inst(memWriteMaskGen_ins_io_inst),
    .io_mask(memWriteMaskGen_ins_io_mask)
  );
  memReadNumGen memReadNumGen_ins ( // @[CtrlUnit.scala 50:33]
    .io_inst(memReadNumGen_ins_io_inst),
    .io_memReadNum(memReadNumGen_ins_io_memReadNum)
  );
  dnpcSrcGen dnpcSrcGen_ins ( // @[CtrlUnit.scala 54:32]
    .io_inst(dnpcSrcGen_ins_io_inst),
    .io_dnpcSrc(dnpcSrcGen_ins_io_dnpcSrc)
  );
  jumpGen jumpGen_ins ( // @[CtrlUnit.scala 58:27]
    .io_inst(jumpGen_ins_io_inst),
    .io_jump(jumpGen_ins_io_jump)
  );
  branchGen branchGen_ins ( // @[CtrlUnit.scala 62:29]
    .io_inst(branchGen_ins_io_inst),
    .io_branch(branchGen_ins_io_branch)
  );
  regEnGen regEnGen_ins ( // @[CtrlUnit.scala 67:28]
    .io_inst(regEnGen_ins_io_inst),
    .io_regEn(regEnGen_ins_io_regEn)
  );
  ResultSrcGen ResultSrcGen_ins ( // @[CtrlUnit.scala 71:32]
    .io_inst(ResultSrcGen_ins_io_inst),
    .io_ResultSrc(ResultSrcGen_ins_io_ResultSrc)
  );
  assign io_CtrlS_AluSrc1 = ALUSrcGen_ins_io_AluSrc1; // @[CtrlUnit.scala 39:20]
  assign io_CtrlS_AluSrc2 = ALUSrcGen_ins_io_AluSrc2; // @[CtrlUnit.scala 40:20]
  assign io_CtrlS_ALUCtrl = ALUCtrl_ins_io_ALUCtrl; // @[CtrlUnit.scala 35:20]
  assign io_CtrlS_memWriteM = memWriteMGen_ins_io_memWriteM; // @[CtrlUnit.scala 44:22]
  assign io_CtrlS_memWriteMask = memWriteMaskGen_ins_io_mask; // @[CtrlUnit.scala 48:25]
  assign io_CtrlS_memReadNum = memReadNumGen_ins_io_memReadNum; // @[CtrlUnit.scala 52:23]
  assign io_CtrlS_dnpcSrc = dnpcSrcGen_ins_io_dnpcSrc; // @[CtrlUnit.scala 56:20]
  assign io_CtrlS_jump = jumpGen_ins_io_jump; // @[CtrlUnit.scala 60:17]
  assign io_CtrlS_branch = branchGen_ins_io_branch; // @[CtrlUnit.scala 64:19]
  assign io_CtrlS_regEn = regEnGen_ins_io_regEn; // @[CtrlUnit.scala 69:18]
  assign io_CtrlS_ResultSrc = ResultSrcGen_ins_io_ResultSrc; // @[CtrlUnit.scala 73:22]
  assign io_CtrlS_fencei = 32'h100f == _io_CtrlS_fencei_T; // @[CtrlUnit.scala 75:30]
  assign ALUCtrl_ins_io_inst = io_inst; // @[CtrlUnit.scala 34:23]
  assign ALUSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 38:25]
  assign memWriteMGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 43:28]
  assign memWriteMaskGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 47:31]
  assign memReadNumGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 51:29]
  assign dnpcSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 55:26]
  assign jumpGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 59:23]
  assign branchGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 63:25]
  assign regEnGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 68:24]
  assign ResultSrcGen_ins_io_inst = io_inst; // @[CtrlUnit.scala 72:28]
endmodule
module csrCtrl(
  input  [31:0] io_inst,
  output        io_CSRCtrlIf_csrrwen,
  output        io_CSRCtrlIf_csrswen,
  output        io_CSRCtrlIf_csrrsien,
  output        io_CSRCtrlIf_csrrcien,
  output        io_CSRCtrlIf_csrrcen,
  output        io_CSRCtrlIf_csrrwien,
  output        io_CSRCtrlIf_ecall,
  output        io_CSRCtrlIf_rfen,
  output        io_CSRCtrlIf_mepc2pc
);
  wire [31:0] _io_CSRCtrlIf_csrrwen_T = io_inst & 32'h707f; // @[csrCtrl.scala 43:35]
  wire  _io_CSRCtrlIf_csrrwen_T_1 = 32'h1073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 43:35]
  wire  _io_CSRCtrlIf_csrswen_T_1 = 32'h2073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 44:35]
  wire  _io_CSRCtrlIf_csrrsien_T_1 = 32'h6073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 45:36]
  wire  _io_CSRCtrlIf_csrrcien_T_1 = 32'h7073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 46:36]
  wire  _io_CSRCtrlIf_csrrcen_T_1 = 32'h3073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 47:35]
  assign io_CSRCtrlIf_csrrwen = 32'h1073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 43:35]
  assign io_CSRCtrlIf_csrswen = 32'h2073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 44:35]
  assign io_CSRCtrlIf_csrrsien = 32'h6073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 45:36]
  assign io_CSRCtrlIf_csrrcien = 32'h7073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 46:36]
  assign io_CSRCtrlIf_csrrcen = 32'h3073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 47:35]
  assign io_CSRCtrlIf_csrrwien = 32'h5073 == _io_CSRCtrlIf_csrrwen_T; // @[csrCtrl.scala 48:36]
  assign io_CSRCtrlIf_ecall = 32'h73 == io_inst; // @[csrCtrl.scala 40:34]
  assign io_CSRCtrlIf_rfen = _io_CSRCtrlIf_csrrwen_T_1 | _io_CSRCtrlIf_csrswen_T_1 | _io_CSRCtrlIf_csrrsien_T_1 |
    _io_CSRCtrlIf_csrrcien_T_1 | _io_CSRCtrlIf_csrrcen_T_1; // @[csrCtrl.scala 50:101]
  assign io_CSRCtrlIf_mepc2pc = 32'h30200073 == io_inst; // @[csrCtrl.scala 52:35]
endmodule
module riscv(
  input          clock,
  input          reset,
  output         io_instIO_valid,
  input          io_instIO_ready,
  input  [63:0]  io_instIO_data_read,
  output [31:0]  io_instIO_addr,
  output         io_dataIO_valid,
  input          io_dataIO_ready,
  input  [63:0]  io_dataIO_data_read,
  output [63:0]  io_dataIO_data_write,
  output         io_dataIO_wen,
  output [31:0]  io_dataIO_addr,
  output [1:0]   io_dataIO_rsize,
  output [7:0]   io_dataIO_mask,
  output         dmaEn_0,
  input          intrTimeCnt_0,
  output         startTimeCnt,
  output [191:0] dmaCtrl,
  input          blockDMA_0,
  output         block2_0,
  output         fencei_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [447:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [191:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[riscv.scala 32:19]
  wire  ifu_reset; // @[riscv.scala 32:19]
  wire [31:0] ifu_io_instIn; // @[riscv.scala 32:19]
  wire [31:0] ifu_io_instOut; // @[riscv.scala 32:19]
  wire [31:0] ifu_io_pc; // @[riscv.scala 32:19]
  wire [31:0] ifu_io_snpc; // @[riscv.scala 32:19]
  wire [31:0] ifu_io_dnpc; // @[riscv.scala 32:19]
  wire  ifu_io_jump; // @[riscv.scala 32:19]
  wire  ifu_intrTimeCnt_0; // @[riscv.scala 32:19]
  wire  ifu_hazardPCBlock_0; // @[riscv.scala 32:19]
  wire  ifu_blockDMA_0; // @[riscv.scala 32:19]
  wire  ifu_block1_0; // @[riscv.scala 32:19]
  wire  ifu_block23_0; // @[riscv.scala 32:19]
  wire  idu_clock; // @[riscv.scala 33:19]
  wire [31:0] idu_io_pc; // @[riscv.scala 33:19]
  wire [31:0] idu_io_inst; // @[riscv.scala 33:19]
  wire  idu_io_regEn; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dataEx_imme; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dataEx_dOut1; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dataEx_dOut2; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dataEx_dIn; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dataEx_rdDout; // @[riscv.scala 33:19]
  wire [4:0] idu_io_rdOut; // @[riscv.scala 33:19]
  wire [4:0] idu_io_rdIn; // @[riscv.scala 33:19]
  wire [4:0] idu_io_rs1; // @[riscv.scala 33:19]
  wire [4:0] idu_io_rs2; // @[riscv.scala 33:19]
  wire [4:0] idu_io_rsWB; // @[riscv.scala 33:19]
  wire [63:0] idu_io_dOutWB; // @[riscv.scala 33:19]
  wire  idu_block1; // @[riscv.scala 33:19]
  wire  idu_block23; // @[riscv.scala 33:19]
  wire  exu_clock; // @[riscv.scala 34:19]
  wire  exu_reset; // @[riscv.scala 34:19]
  wire [1:0] exu_io_AluSrc1; // @[riscv.scala 34:19]
  wire [1:0] exu_io_AluSrc2; // @[riscv.scala 34:19]
  wire [4:0] exu_io_ALUCtrl; // @[riscv.scala 34:19]
  wire  exu_io_dnpcSrc; // @[riscv.scala 34:19]
  wire [1:0] exu_io_ResultSrc; // @[riscv.scala 34:19]
  wire [2:0] exu_io_memReadNum; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataId_imme; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataId_dOut1; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataId_dOut2; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataId_dIn; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataId_rdDout; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataOut_ALUResOut; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataOut_wdata; // @[riscv.scala 34:19]
  wire [63:0] exu_io_dataOut_rdata; // @[riscv.scala 34:19]
  wire  exu_io_brTake; // @[riscv.scala 34:19]
  wire [31:0] exu_io_pc; // @[riscv.scala 34:19]
  wire [31:0] exu_io_snpc; // @[riscv.scala 34:19]
  wire [31:0] exu_io_dnpc; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrrwen; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrswen; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrrsien; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrrcien; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrrcen; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_csrrwien; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_ecall; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_rfen; // @[riscv.scala 34:19]
  wire  exu_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 34:19]
  wire [4:0] exu_io_uimm; // @[riscv.scala 34:19]
  wire [63:0] exu_io_aluResIn; // @[riscv.scala 34:19]
  wire [1:0] exu_io_forwardA; // @[riscv.scala 34:19]
  wire [1:0] exu_io_forwardB; // @[riscv.scala 34:19]
  wire [1:0] exu_io_forwardC; // @[riscv.scala 34:19]
  wire [63:0] exu_io_aluRes1; // @[riscv.scala 34:19]
  wire [63:0] exu_io_aluRes3; // @[riscv.scala 34:19]
  wire  exu_intrTimeCnt_0; // @[riscv.scala 34:19]
  wire  exu_startTimeCnt; // @[riscv.scala 34:19]
  wire [191:0] exu_dmaCtrl_0; // @[riscv.scala 34:19]
  wire  exu_blockDMA; // @[riscv.scala 34:19]
  wire  exu_block1; // @[riscv.scala 34:19]
  wire  exu_block23; // @[riscv.scala 34:19]
  wire  hazardu_io_regEnEXMEM; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rdEXMEM; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rs1IDEX; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rs2IDEX; // @[riscv.scala 35:23]
  wire  hazardu_io_regEnMEMWB; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rdMEMWB; // @[riscv.scala 35:23]
  wire  hazardu_io_regEnWBEND; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rdWBEND; // @[riscv.scala 35:23]
  wire [1:0] hazardu_io_forwardA; // @[riscv.scala 35:23]
  wire [1:0] hazardu_io_forwardB; // @[riscv.scala 35:23]
  wire [1:0] hazardu_io_forwardC; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rs1IFID; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rs2IFID; // @[riscv.scala 35:23]
  wire [4:0] hazardu_io_rdIDEX; // @[riscv.scala 35:23]
  wire [1:0] hazardu_io_resSrc; // @[riscv.scala 35:23]
  wire  hazardu_io_loadHazard; // @[riscv.scala 35:23]
  wire  preBranchIns_clock; // @[riscv.scala 36:28]
  wire  preBranchIns_reset; // @[riscv.scala 36:28]
  wire  preBranchIns_io_exjump; // @[riscv.scala 36:28]
  wire [31:0] preBranchIns_io_ifpc; // @[riscv.scala 36:28]
  wire [31:0] preBranchIns_io_expc; // @[riscv.scala 36:28]
  wire [31:0] preBranchIns_io_exdpc; // @[riscv.scala 36:28]
  wire [31:0] preBranchIns_io_ifdnpc; // @[riscv.scala 36:28]
  wire  preBranchIns_io_ifjump; // @[riscv.scala 36:28]
  wire  preBranchIns_block1_0; // @[riscv.scala 36:28]
  wire  preBranchIns_block23_0; // @[riscv.scala 36:28]
  wire [31:0] memVGenInst_io_inst; // @[riscv.scala 60:28]
  wire  memVGenInst_io_valid; // @[riscv.scala 60:28]
  wire [31:0] ctrl_io_inst; // @[riscv.scala 65:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc1; // @[riscv.scala 65:20]
  wire [1:0] ctrl_io_CtrlS_AluSrc2; // @[riscv.scala 65:20]
  wire [4:0] ctrl_io_CtrlS_ALUCtrl; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_memWriteM; // @[riscv.scala 65:20]
  wire [7:0] ctrl_io_CtrlS_memWriteMask; // @[riscv.scala 65:20]
  wire [2:0] ctrl_io_CtrlS_memReadNum; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_dnpcSrc; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_jump; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_branch; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_regEn; // @[riscv.scala 65:20]
  wire [1:0] ctrl_io_CtrlS_ResultSrc; // @[riscv.scala 65:20]
  wire  ctrl_io_CtrlS_fencei; // @[riscv.scala 65:20]
  wire [31:0] csrCtrl_io_inst; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwen; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrswen; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrsien; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcien; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrcen; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_csrrwien; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_ecall; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_rfen; // @[riscv.scala 66:23]
  wire  csrCtrl_io_CSRCtrlIf_mepc2pc; // @[riscv.scala 66:23]
  wire  difftest_v; // @[riscv.scala 384:24]
  wire  intrins_intr; // @[riscv.scala 390:23]
  wire  Ebpro_block; // @[riscv.scala 396:21]
  wire [31:0] Ebpro_inst; // @[riscv.scala 396:21]
  wire  skipinst_v; // @[riscv.scala 400:24]
  wire  block1_0 = exu_block1;
  wire  _io_instIO_valid_T = ~block1_0; // @[riscv.scala 53:32]
  wire  _io_instIO_valid_T_2 = ~blockDMA_0; // @[riscv.scala 53:43]
  wire  _block2_T_1 = ~io_instIO_ready; // @[riscv.scala 57:23]
  wire  block2 = ~io_instIO_ready; // @[riscv.scala 57:23]
  reg [248:0] pipEX2MEMReg; // @[Reg.scala 27:20]
  wire  pipEX2MEMWire_valid = pipEX2MEMReg[47]; // @[riscv.scala 253:44]
  wire  block3 = pipEX2MEMWire_valid & ~io_dataIO_ready; // @[riscv.scala 268:33]
  wire  block23 = _block2_T_1 | block3; // @[riscv.scala 273:21]
  wire  pipBlock = block1_0 | block23 | blockDMA_0; // @[riscv.scala 376:32]
  wire  _T = ~pipBlock; // @[riscv.scala 86:30]
  reg [430:0] pipID2ExReg; // @[Reg.scala 27:20]
  wire  pipID2ExWire_branch = pipID2ExReg[48]; // @[riscv.scala 163:41]
  wire  pipID2ExWire_jump = pipID2ExReg[49]; // @[riscv.scala 163:41]
  reg [8:0] pipCSRReg; // @[Reg.scala 27:20]
  wire  pipCSRRegWire_mepc2pc = pipCSRReg[0]; // @[riscv.scala 210:41]
  wire  pipCSRRegWire_ecall = pipCSRReg[2]; // @[riscv.scala 210:41]
  wire  dnpcTakenWithoutPreB = pipID2ExWire_branch & exu_io_brTake | pipID2ExWire_jump | pipCSRRegWire_mepc2pc |
    pipCSRRegWire_ecall; // @[riscv.scala 330:115]
  wire  pipID2ExWire_ifjump = pipID2ExReg[33]; // @[riscv.scala 163:41]
  wire  jump1 = ~dnpcTakenWithoutPreB & pipID2ExWire_ifjump; // @[riscv.scala 331:37]
  wire [31:0] pipID2ExWire_ifdnpc = pipID2ExReg[32:1]; // @[riscv.scala 163:41]
  wire  jump2 = dnpcTakenWithoutPreB & (exu_io_dnpc != pipID2ExWire_ifdnpc | ~pipID2ExWire_ifjump); // @[riscv.scala 332:36]
  wire [31:0] pipID2ExWire_pc = pipID2ExReg[141:110]; // @[riscv.scala 163:41]
  wire  _pipFlashWire_T_2 = intrTimeCnt_0 & pipID2ExWire_pc != 32'h0; // @[riscv.scala 333:50]
  wire  pipID2ExWire_fencei = pipID2ExReg[34]; // @[riscv.scala 163:41]
  wire  pipFlashWire = jump1 | jump2 | intrTimeCnt_0 & pipID2ExWire_pc != 32'h0 | pipID2ExWire_fencei; // @[riscv.scala 333:78]
  wire  _T_3 = pipFlashWire & ~pipBlock | reset; // @[riscv.scala 86:40]
  wire  pipIF2IDReg_hi_hi_hi = ifu_io_pc != 32'h0; // @[riscv.scala 88:16]
  wire [129:0] _pipIF2IDReg_T = {pipIF2IDReg_hi_hi_hi,ifu_io_instOut,ifu_io_pc,ifu_io_snpc,preBranchIns_io_ifjump,
    preBranchIns_io_ifdnpc}; // @[Cat.scala 30:58]
  wire  _pipIF2IDReg_T_2 = ~(pipBlock | hazardu_io_loadHazard); // @[riscv.scala 94:13]
  reg [129:0] pipIF2IDReg; // @[Reg.scala 27:20]
  wire [31:0] pipIF2IDWire_ifdnpc = pipIF2IDReg[31:0]; // @[riscv.scala 96:41]
  wire  pipIF2IDWire_ifjump = pipIF2IDReg[32]; // @[riscv.scala 96:41]
  wire [31:0] pipIF2IDWire_snpc = pipIF2IDReg[64:33]; // @[riscv.scala 96:41]
  wire [31:0] pipIF2IDWire_pc = pipIF2IDReg[96:65]; // @[riscv.scala 96:41]
  wire [31:0] pipIF2IDWire_inst = pipIF2IDReg[128:97]; // @[riscv.scala 96:41]
  wire  pipIF2IDWire_cmd = pipIF2IDReg[129]; // @[riscv.scala 96:41]
  wire  _T_8 = (pipFlashWire | hazardu_io_loadHazard) & _T | reset; // @[riscv.scala 131:67]
  wire [31:0] _pipID2ExReg_T = pipIF2IDWire_inst & 32'hfe00707f; // @[riscv.scala 159:25]
  wire  pipID2ExReg_lo_lo_lo_lo = 32'hc00607b == _pipID2ExReg_T; // @[riscv.scala 159:25]
  wire [44:0] pipID2ExReg_lo_lo = {idu_io_rs1,idu_io_rs2,ctrl_io_CtrlS_fencei,pipIF2IDWire_ifjump,pipIF2IDWire_ifdnpc,
    pipID2ExReg_lo_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [59:0] pipID2ExReg_lo = {ctrl_io_CtrlS_memWriteMask,ctrl_io_CtrlS_memWriteM,ctrl_io_CtrlS_dnpcSrc,
    ctrl_io_CtrlS_jump,ctrl_io_CtrlS_branch,ctrl_io_CtrlS_regEn,ctrl_io_CtrlS_ResultSrc,pipID2ExReg_lo_lo}; // @[Cat.scala 30:58]
  wire [49:0] pipID2ExReg_hi_lo = {pipIF2IDWire_snpc,idu_io_rdOut,ctrl_io_CtrlS_ALUCtrl,ctrl_io_CtrlS_AluSrc1,
    ctrl_io_CtrlS_AluSrc2,ctrl_io_CtrlS_memReadNum,memVGenInst_io_valid}; // @[Cat.scala 30:58]
  wire [430:0] _pipID2ExReg_T_1 = {pipIF2IDWire_cmd,pipIF2IDWire_inst,idu_io_dataEx_imme,idu_io_dataEx_dOut1,
    idu_io_dataEx_dOut2,idu_io_dataEx_rdDout,pipIF2IDWire_pc,pipID2ExReg_hi_lo,pipID2ExReg_lo}; // @[Cat.scala 30:58]
  wire  pipID2ExWire_dma = pipID2ExReg[0]; // @[riscv.scala 163:41]
  wire [1:0] pipID2ExWire_resultSrc = pipID2ExReg[46:45]; // @[riscv.scala 163:41]
  wire  pipID2ExWire_regEn = pipID2ExReg[47]; // @[riscv.scala 163:41]
  wire  pipID2ExWire_memWriteM = pipID2ExReg[51]; // @[riscv.scala 163:41]
  wire [7:0] pipID2ExWire_mask = pipID2ExReg[59:52]; // @[riscv.scala 163:41]
  wire  pipID2ExWire_valid = pipID2ExReg[60]; // @[riscv.scala 163:41]
  wire [2:0] pipID2ExWire_memReadNum = pipID2ExReg[63:61]; // @[riscv.scala 163:41]
  wire [4:0] pipID2ExWire_rd = pipID2ExReg[77:73]; // @[riscv.scala 163:41]
  wire [31:0] pipID2ExWire_snpc = pipID2ExReg[109:78]; // @[riscv.scala 163:41]
  wire [31:0] pipID2ExWire_inst = pipID2ExReg[429:398]; // @[riscv.scala 163:41]
  wire  pipID2ExWire_cmd = pipID2ExReg[430]; // @[riscv.scala 163:41]
  wire [8:0] _pipCSRReg_T = {csrCtrl_io_CSRCtrlIf_csrrwen,csrCtrl_io_CSRCtrlIf_csrswen,csrCtrl_io_CSRCtrlIf_csrrsien,
    csrCtrl_io_CSRCtrlIf_csrrcien,csrCtrl_io_CSRCtrlIf_csrrcen,csrCtrl_io_CSRCtrlIf_csrrwien,csrCtrl_io_CSRCtrlIf_ecall,
    csrCtrl_io_CSRCtrlIf_rfen,csrCtrl_io_CSRCtrlIf_mepc2pc}; // @[Cat.scala 30:58]
  wire  pipCSRRegWire_rfen = pipCSRReg[1]; // @[riscv.scala 210:41]
  wire  pipEX2MEMReg_lo_hi_lo_hi = pipID2ExWire_regEn | pipCSRRegWire_rfen; // @[riscv.scala 246:21]
  wire  _pipID2ExWire_WIRE_dma = pipID2ExWire_dma; // @[riscv.scala 163:41]
  wire [46:0] pipEX2MEMReg_lo = {pipID2ExWire_mask,pipID2ExWire_memWriteM,pipEX2MEMReg_lo_hi_lo_hi,
    pipID2ExWire_resultSrc,pipID2ExWire_pc,pipID2ExWire_fencei,_pipFlashWire_T_2,pipID2ExWire_dma}; // @[Cat.scala 30:58]
  wire [248:0] _pipEX2MEMReg_T_3 = {pipID2ExWire_cmd,pipID2ExWire_inst,exu_io_dataOut_ALUResOut,exu_io_dataOut_wdata,
    pipID2ExWire_snpc,pipID2ExWire_rd,pipID2ExWire_memReadNum,pipID2ExWire_valid,pipEX2MEMReg_lo}; // @[Cat.scala 30:58]
  wire  pipEX2MEMWire_skip = pipEX2MEMReg[0]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_intr = pipEX2MEMReg[1]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_fencei = pipEX2MEMReg[2]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_pc = pipEX2MEMReg[34:3]; // @[riscv.scala 253:44]
  wire [1:0] pipEX2MEMWire_ResultSrc = pipEX2MEMReg[36:35]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_regEn = pipEX2MEMReg[37]; // @[riscv.scala 253:44]
  wire [7:0] pipEX2MEMWire_mask = pipEX2MEMReg[46:39]; // @[riscv.scala 253:44]
  wire [2:0] pipEX2MEMWire_memReadNum = pipEX2MEMReg[50:48]; // @[riscv.scala 253:44]
  wire [4:0] pipEX2MEMWire_rd = pipEX2MEMReg[55:51]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_snpc = pipEX2MEMReg[87:56]; // @[riscv.scala 253:44]
  wire [63:0] pipEX2MEMWire_writeDataM = pipEX2MEMReg[151:88]; // @[riscv.scala 253:44]
  wire [63:0] pipEX2MEMWire_ALURes = pipEX2MEMReg[215:152]; // @[riscv.scala 253:44]
  wire [31:0] pipEX2MEMWire_inst = pipEX2MEMReg[247:216]; // @[riscv.scala 253:44]
  wire  pipEX2MEMWire_cmd = pipEX2MEMReg[248]; // @[riscv.scala 253:44]
  wire [14:0] _GEN_7 = {{7'd0}, pipEX2MEMWire_mask}; // @[riscv.scala 256:40]
  wire [14:0] _io_dataIO_mask_T_1 = _GEN_7 << pipEX2MEMWire_ALURes[2:0]; // @[riscv.scala 256:40]
  wire [6:0] _io_dataIO_data_write_T_1 = pipEX2MEMWire_ALURes[2:0] * 4'h8; // @[riscv.scala 261:78]
  wire [190:0] _GEN_8 = {{127'd0}, pipEX2MEMWire_writeDataM}; // @[riscv.scala 261:50]
  wire [190:0] _io_dataIO_data_write_T_2 = _GEN_8 << _io_dataIO_data_write_T_1; // @[riscv.scala 261:50]
  wire  skip = pipEX2MEMWire_valid & (pipEX2MEMWire_ALURes < 64'h80000000 | pipEX2MEMWire_ALURes > 64'h8fffffff) |
    pipEX2MEMWire_fencei; // @[riscv.scala 265:109]
  wire  jud = pipEX2MEMWire_pc == 32'h0; // @[riscv.scala 278:29]
  wire  pipMEM2WBReg_lo_lo_lo = skip | pipEX2MEMWire_skip; // @[riscv.scala 291:10]
  reg [173:0] pipMEM2WBReg; // @[Reg.scala 27:20]
  wire [31:0] pipMEM2WBWire_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 293:44]
  wire [31:0] _lo_T_1 = pipMEM2WBWire_pc + 32'h4; // @[riscv.scala 294:42]
  wire [31:0] npcsend = jud ? _lo_T_1 : pipEX2MEMWire_pc; // @[riscv.scala 294:17]
  wire [36:0] pipMEM2WBReg_lo = {pipEX2MEMWire_regEn,pipEX2MEMWire_ResultSrc,npcsend,pipEX2MEMWire_intr,
    pipMEM2WBReg_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [173:0] _pipMEM2WBReg_T = {pipEX2MEMWire_cmd,pipEX2MEMWire_inst,pipEX2MEMWire_ALURes,pipEX2MEMWire_rd,
    pipEX2MEMWire_snpc,pipEX2MEMWire_memReadNum,pipMEM2WBReg_lo}; // @[Cat.scala 30:58]
  wire  pipMEM2WBWire_intr = pipMEM2WBReg[1]; // @[riscv.scala 293:44]
  wire  pipMEM2WBWire_regEn = pipMEM2WBReg[36]; // @[riscv.scala 293:44]
  wire [4:0] pipMEM2WBWire_rd = pipMEM2WBReg[76:72]; // @[riscv.scala 293:44]
  wire [63:0] pipMEM2WBWire_ALURes = pipMEM2WBReg[140:77]; // @[riscv.scala 293:44]
  wire [31:0] pipMEM2WBWire_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 293:44]
  wire  pipMEM2WBWire_cmd = pipMEM2WBReg[173]; // @[riscv.scala 293:44]
  reg [63:0] exu_io_dataOut_rdata_r; // @[Reg.scala 27:20]
  wire [6:0] _exu_io_dataOut_rdata_T_2 = pipMEM2WBWire_ALURes[2:0] * 4'h8; // @[riscv.scala 302:100]
  wire [69:0] _pipWB2ENDWire_T = {pipMEM2WBWire_rd,pipMEM2WBWire_regEn,pipMEM2WBWire_inst,pipMEM2WBWire_pc}; // @[Cat.scala 30:58]
  reg [69:0] pipWB2ENDWire_r; // @[Reg.scala 27:20]
  wire [31:0] _ifu_io_dnpc_T_2 = jump2 ? exu_io_dnpc : preBranchIns_io_ifdnpc; // @[riscv.scala 345:12]
  wire [31:0] _ifu_io_dnpc_T_3 = jump1 ? pipID2ExWire_snpc : _ifu_io_dnpc_T_2; // @[riscv.scala 342:10]
  wire [31:0] _ifu_io_dnpc_T_4 = pipID2ExWire_fencei ? pipID2ExWire_snpc : _ifu_io_dnpc_T_3; // @[riscv.scala 339:8]
  wire  hazardPCBlock = hazardu_io_loadHazard; // @[riscv.scala 372:27 riscv.scala 373:17]
  wire  dmaEn = pipID2ExWire_dma; // @[riscv.scala 163:41]
  wire  fencei = pipID2ExWire_fencei & ~intrTimeCnt_0 & _T; // @[riscv.scala 379:49]
  iFetch ifu ( // @[riscv.scala 32:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_instIn(ifu_io_instIn),
    .io_instOut(ifu_io_instOut),
    .io_pc(ifu_io_pc),
    .io_snpc(ifu_io_snpc),
    .io_dnpc(ifu_io_dnpc),
    .io_jump(ifu_io_jump),
    .intrTimeCnt_0(ifu_intrTimeCnt_0),
    .hazardPCBlock_0(ifu_hazardPCBlock_0),
    .blockDMA_0(ifu_blockDMA_0),
    .block1_0(ifu_block1_0),
    .block23_0(ifu_block23_0)
  );
  iDecode idu ( // @[riscv.scala 33:19]
    .clock(idu_clock),
    .io_pc(idu_io_pc),
    .io_inst(idu_io_inst),
    .io_regEn(idu_io_regEn),
    .io_dataEx_imme(idu_io_dataEx_imme),
    .io_dataEx_dOut1(idu_io_dataEx_dOut1),
    .io_dataEx_dOut2(idu_io_dataEx_dOut2),
    .io_dataEx_dIn(idu_io_dataEx_dIn),
    .io_dataEx_rdDout(idu_io_dataEx_rdDout),
    .io_rdOut(idu_io_rdOut),
    .io_rdIn(idu_io_rdIn),
    .io_rs1(idu_io_rs1),
    .io_rs2(idu_io_rs2),
    .io_rsWB(idu_io_rsWB),
    .io_dOutWB(idu_io_dOutWB),
    .block1(idu_block1),
    .block23(idu_block23)
  );
  execute exu ( // @[riscv.scala 34:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_AluSrc1(exu_io_AluSrc1),
    .io_AluSrc2(exu_io_AluSrc2),
    .io_ALUCtrl(exu_io_ALUCtrl),
    .io_dnpcSrc(exu_io_dnpcSrc),
    .io_ResultSrc(exu_io_ResultSrc),
    .io_memReadNum(exu_io_memReadNum),
    .io_dataId_imme(exu_io_dataId_imme),
    .io_dataId_dOut1(exu_io_dataId_dOut1),
    .io_dataId_dOut2(exu_io_dataId_dOut2),
    .io_dataId_dIn(exu_io_dataId_dIn),
    .io_dataId_rdDout(exu_io_dataId_rdDout),
    .io_dataOut_ALUResOut(exu_io_dataOut_ALUResOut),
    .io_dataOut_wdata(exu_io_dataOut_wdata),
    .io_dataOut_rdata(exu_io_dataOut_rdata),
    .io_brTake(exu_io_brTake),
    .io_pc(exu_io_pc),
    .io_snpc(exu_io_snpc),
    .io_dnpc(exu_io_dnpc),
    .io_CSRCtrlIf_csrrwen(exu_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(exu_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(exu_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(exu_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(exu_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(exu_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(exu_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(exu_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(exu_io_CSRCtrlIf_mepc2pc),
    .io_uimm(exu_io_uimm),
    .io_aluResIn(exu_io_aluResIn),
    .io_forwardA(exu_io_forwardA),
    .io_forwardB(exu_io_forwardB),
    .io_forwardC(exu_io_forwardC),
    .io_aluRes1(exu_io_aluRes1),
    .io_aluRes3(exu_io_aluRes3),
    .intrTimeCnt_0(exu_intrTimeCnt_0),
    .startTimeCnt(exu_startTimeCnt),
    .dmaCtrl_0(exu_dmaCtrl_0),
    .blockDMA(exu_blockDMA),
    .block1(exu_block1),
    .block23(exu_block23)
  );
  hazard hazardu ( // @[riscv.scala 35:23]
    .io_regEnEXMEM(hazardu_io_regEnEXMEM),
    .io_rdEXMEM(hazardu_io_rdEXMEM),
    .io_rs1IDEX(hazardu_io_rs1IDEX),
    .io_rs2IDEX(hazardu_io_rs2IDEX),
    .io_regEnMEMWB(hazardu_io_regEnMEMWB),
    .io_rdMEMWB(hazardu_io_rdMEMWB),
    .io_regEnWBEND(hazardu_io_regEnWBEND),
    .io_rdWBEND(hazardu_io_rdWBEND),
    .io_forwardA(hazardu_io_forwardA),
    .io_forwardB(hazardu_io_forwardB),
    .io_forwardC(hazardu_io_forwardC),
    .io_rs1IFID(hazardu_io_rs1IFID),
    .io_rs2IFID(hazardu_io_rs2IFID),
    .io_rdIDEX(hazardu_io_rdIDEX),
    .io_resSrc(hazardu_io_resSrc),
    .io_loadHazard(hazardu_io_loadHazard)
  );
  preBranch preBranchIns ( // @[riscv.scala 36:28]
    .clock(preBranchIns_clock),
    .reset(preBranchIns_reset),
    .io_exjump(preBranchIns_io_exjump),
    .io_ifpc(preBranchIns_io_ifpc),
    .io_expc(preBranchIns_io_expc),
    .io_exdpc(preBranchIns_io_exdpc),
    .io_ifdnpc(preBranchIns_io_ifdnpc),
    .io_ifjump(preBranchIns_io_ifjump),
    .block1_0(preBranchIns_block1_0),
    .block23_0(preBranchIns_block23_0)
  );
  memVGen memVGenInst ( // @[riscv.scala 60:28]
    .io_inst(memVGenInst_io_inst),
    .io_valid(memVGenInst_io_valid)
  );
  CtrlUnit ctrl ( // @[riscv.scala 65:20]
    .io_inst(ctrl_io_inst),
    .io_CtrlS_AluSrc1(ctrl_io_CtrlS_AluSrc1),
    .io_CtrlS_AluSrc2(ctrl_io_CtrlS_AluSrc2),
    .io_CtrlS_ALUCtrl(ctrl_io_CtrlS_ALUCtrl),
    .io_CtrlS_memWriteM(ctrl_io_CtrlS_memWriteM),
    .io_CtrlS_memWriteMask(ctrl_io_CtrlS_memWriteMask),
    .io_CtrlS_memReadNum(ctrl_io_CtrlS_memReadNum),
    .io_CtrlS_dnpcSrc(ctrl_io_CtrlS_dnpcSrc),
    .io_CtrlS_jump(ctrl_io_CtrlS_jump),
    .io_CtrlS_branch(ctrl_io_CtrlS_branch),
    .io_CtrlS_regEn(ctrl_io_CtrlS_regEn),
    .io_CtrlS_ResultSrc(ctrl_io_CtrlS_ResultSrc),
    .io_CtrlS_fencei(ctrl_io_CtrlS_fencei)
  );
  csrCtrl csrCtrl ( // @[riscv.scala 66:23]
    .io_inst(csrCtrl_io_inst),
    .io_CSRCtrlIf_csrrwen(csrCtrl_io_CSRCtrlIf_csrrwen),
    .io_CSRCtrlIf_csrswen(csrCtrl_io_CSRCtrlIf_csrswen),
    .io_CSRCtrlIf_csrrsien(csrCtrl_io_CSRCtrlIf_csrrsien),
    .io_CSRCtrlIf_csrrcien(csrCtrl_io_CSRCtrlIf_csrrcien),
    .io_CSRCtrlIf_csrrcen(csrCtrl_io_CSRCtrlIf_csrrcen),
    .io_CSRCtrlIf_csrrwien(csrCtrl_io_CSRCtrlIf_csrrwien),
    .io_CSRCtrlIf_ecall(csrCtrl_io_CSRCtrlIf_ecall),
    .io_CSRCtrlIf_rfen(csrCtrl_io_CSRCtrlIf_rfen),
    .io_CSRCtrlIf_mepc2pc(csrCtrl_io_CSRCtrlIf_mepc2pc)
  );
  difftest difftest ( // @[riscv.scala 384:24]
    .v(difftest_v)
  );
  intr intrins ( // @[riscv.scala 390:23]
    .intr(intrins_intr)
  );
  ebProbe Ebpro ( // @[riscv.scala 396:21]
    .block(Ebpro_block),
    .inst(Ebpro_inst)
  );
  skip skipinst ( // @[riscv.scala 400:24]
    .v(skipinst_v)
  );
  assign io_instIO_valid = ~block1_0 & ~blockDMA_0; // @[riscv.scala 53:40]
  assign io_instIO_addr = ifu_io_pc; // @[riscv.scala 79:18]
  assign io_dataIO_valid = pipEX2MEMWire_valid & _io_instIO_valid_T & _io_instIO_valid_T_2; // @[riscv.scala 262:53]
  assign io_dataIO_data_write = _io_dataIO_data_write_T_2[63:0]; // @[riscv.scala 261:23]
  assign io_dataIO_wen = pipEX2MEMReg[38]; // @[riscv.scala 253:44]
  assign io_dataIO_addr = pipEX2MEMWire_ALURes[31:0]; // @[riscv.scala 259:18]
  assign io_dataIO_rsize = pipEX2MEMWire_memReadNum[1:0]; // @[riscv.scala 260:46]
  assign io_dataIO_mask = _io_dataIO_mask_T_1[7:0]; // @[riscv.scala 256:18]
  assign dmaEn_0 = _pipID2ExWire_WIRE_dma;
  assign startTimeCnt = exu_startTimeCnt;
  assign dmaCtrl = exu_dmaCtrl_0;
  assign block2_0 = _block2_T_1;
  assign fencei_0 = fencei;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_instIn = ifu_io_pc[2] ? io_instIO_data_read[63:32] : io_instIO_data_read[31:0]; // @[riscv.scala 78:23]
  assign ifu_io_dnpc = _pipFlashWire_T_2 ? exu_io_dnpc : _ifu_io_dnpc_T_4; // @[riscv.scala 336:21]
  assign ifu_io_jump = pipFlashWire | preBranchIns_io_ifjump; // @[riscv.scala 335:100]
  assign ifu_intrTimeCnt_0 = intrTimeCnt_0;
  assign ifu_hazardPCBlock_0 = hazardPCBlock;
  assign ifu_blockDMA_0 = blockDMA_0;
  assign ifu_block1_0 = exu_block1;
  assign ifu_block23_0 = block23;
  assign idu_clock = clock;
  assign idu_io_pc = pipMEM2WBReg[33:2]; // @[riscv.scala 293:44]
  assign idu_io_inst = pipIF2IDReg[128:97]; // @[riscv.scala 96:41]
  assign idu_io_regEn = pipMEM2WBReg[36]; // @[riscv.scala 293:44]
  assign idu_io_dataEx_dIn = exu_io_dataId_dIn; // @[riscv.scala 303:21]
  assign idu_io_rdIn = pipMEM2WBReg[76:72]; // @[riscv.scala 293:44]
  assign idu_io_rsWB = pipWB2ENDWire_r[69:65]; // @[riscv.scala 324:13]
  assign idu_block1 = exu_block1;
  assign idu_block23 = block23;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_AluSrc1 = pipID2ExReg[67:66]; // @[riscv.scala 163:41]
  assign exu_io_AluSrc2 = pipID2ExReg[65:64]; // @[riscv.scala 163:41]
  assign exu_io_ALUCtrl = pipID2ExReg[72:68]; // @[riscv.scala 163:41]
  assign exu_io_dnpcSrc = pipID2ExReg[50]; // @[riscv.scala 163:41]
  assign exu_io_ResultSrc = pipMEM2WBReg[35:34]; // @[riscv.scala 293:44]
  assign exu_io_memReadNum = pipMEM2WBReg[39:37]; // @[riscv.scala 293:44]
  assign exu_io_dataId_imme = pipID2ExReg[397:334]; // @[riscv.scala 163:41]
  assign exu_io_dataId_dOut1 = pipID2ExReg[333:270]; // @[riscv.scala 163:41]
  assign exu_io_dataId_dOut2 = pipID2ExReg[269:206]; // @[riscv.scala 163:41]
  assign exu_io_dataId_rdDout = pipID2ExReg[205:142]; // @[riscv.scala 163:41]
  assign exu_io_dataOut_rdata = exu_io_dataOut_rdata_r >> _exu_io_dataOut_rdata_T_2; // @[riscv.scala 302:73]
  assign exu_io_pc = pipID2ExReg[141:110]; // @[riscv.scala 163:41]
  assign exu_io_snpc = pipMEM2WBReg[71:40]; // @[riscv.scala 293:44]
  assign exu_io_CSRCtrlIf_csrrwen = pipCSRReg[8]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_csrswen = pipCSRReg[7]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_csrrsien = pipCSRReg[6]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_csrrcien = pipCSRReg[5]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_csrrcen = pipCSRReg[4]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_csrrwien = pipCSRReg[3]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_ecall = pipCSRReg[2]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_rfen = pipCSRReg[1]; // @[riscv.scala 210:41]
  assign exu_io_CSRCtrlIf_mepc2pc = pipCSRReg[0]; // @[riscv.scala 210:41]
  assign exu_io_uimm = pipID2ExReg[44:40]; // @[riscv.scala 163:41]
  assign exu_io_aluResIn = pipMEM2WBReg[140:77]; // @[riscv.scala 293:44]
  assign exu_io_forwardA = hazardu_io_forwardA; // @[riscv.scala 362:19]
  assign exu_io_forwardB = hazardu_io_forwardB; // @[riscv.scala 363:19]
  assign exu_io_forwardC = hazardu_io_forwardC; // @[riscv.scala 364:19]
  assign exu_io_aluRes1 = pipEX2MEMWire_ResultSrc == 2'h0 ? pipEX2MEMWire_ALURes : {{32'd0}, pipEX2MEMWire_snpc}; // @[riscv.scala 263:24]
  assign exu_io_aluRes3 = idu_io_dOutWB; // @[riscv.scala 326:18]
  assign exu_intrTimeCnt_0 = intrTimeCnt_0;
  assign exu_blockDMA = blockDMA_0;
  assign exu_block23 = block23;
  assign hazardu_io_regEnEXMEM = pipEX2MEMReg[37]; // @[riscv.scala 253:44]
  assign hazardu_io_rdEXMEM = pipEX2MEMReg[55:51]; // @[riscv.scala 253:44]
  assign hazardu_io_rs1IDEX = pipID2ExReg[44:40]; // @[riscv.scala 163:41]
  assign hazardu_io_rs2IDEX = pipID2ExReg[39:35]; // @[riscv.scala 163:41]
  assign hazardu_io_regEnMEMWB = pipMEM2WBReg[36]; // @[riscv.scala 293:44]
  assign hazardu_io_rdMEMWB = pipMEM2WBReg[76:72]; // @[riscv.scala 293:44]
  assign hazardu_io_regEnWBEND = pipWB2ENDWire_r[64]; // @[riscv.scala 324:13]
  assign hazardu_io_rdWBEND = pipWB2ENDWire_r[69:65]; // @[riscv.scala 324:13]
  assign hazardu_io_rs1IFID = idu_io_rs1; // @[riscv.scala 367:22]
  assign hazardu_io_rs2IFID = idu_io_rs2; // @[riscv.scala 368:22]
  assign hazardu_io_rdIDEX = pipID2ExReg[77:73]; // @[riscv.scala 163:41]
  assign hazardu_io_resSrc = pipID2ExReg[46:45]; // @[riscv.scala 163:41]
  assign preBranchIns_clock = clock;
  assign preBranchIns_reset = reset;
  assign preBranchIns_io_exjump = pipID2ExWire_branch & exu_io_brTake | pipID2ExWire_jump | pipCSRRegWire_mepc2pc |
    pipCSRRegWire_ecall; // @[riscv.scala 330:115]
  assign preBranchIns_io_ifpc = ifu_io_pc; // @[riscv.scala 404:24]
  assign preBranchIns_io_expc = pipID2ExReg[141:110]; // @[riscv.scala 163:41]
  assign preBranchIns_io_exdpc = exu_io_dnpc; // @[riscv.scala 407:25]
  assign preBranchIns_block1_0 = exu_block1;
  assign preBranchIns_block23_0 = block23;
  assign memVGenInst_io_inst = pipIF2IDReg[128:97]; // @[riscv.scala 96:41]
  assign ctrl_io_inst = pipIF2IDReg[128:97]; // @[riscv.scala 96:41]
  assign csrCtrl_io_inst = pipIF2IDReg[128:97]; // @[riscv.scala 96:41]
  assign difftest_v = pipMEM2WBWire_cmd & _T; // @[riscv.scala 385:38]
  assign intrins_intr = pipMEM2WBWire_intr & _T; // @[riscv.scala 391:41]
  assign Ebpro_block = block1_0 | block23 | blockDMA_0; // @[riscv.scala 376:32]
  assign Ebpro_inst = pipMEM2WBReg[172:141]; // @[riscv.scala 293:44]
  assign skipinst_v = pipMEM2WBReg[0]; // @[riscv.scala 293:44]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      pipEX2MEMReg <= 249'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      if (_pipFlashWire_T_2) begin // @[riscv.scala 232:35]
        pipEX2MEMReg <= 249'h1;
      end else begin
        pipEX2MEMReg <= _pipEX2MEMReg_T_3;
      end
    end
    if (_T_8) begin // @[Reg.scala 27:20]
      pipID2ExReg <= 431'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      pipID2ExReg <= _pipID2ExReg_T_1; // @[Reg.scala 28:23]
    end
    if (_T_8) begin // @[Reg.scala 27:20]
      pipCSRReg <= 9'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      pipCSRReg <= _pipCSRReg_T; // @[Reg.scala 28:23]
    end
    if (_T_3) begin // @[Reg.scala 27:20]
      pipIF2IDReg <= 130'h0; // @[Reg.scala 27:20]
    end else if (_pipIF2IDReg_T_2) begin // @[Reg.scala 28:19]
      pipIF2IDReg <= _pipIF2IDReg_T; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pipMEM2WBReg <= 174'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      pipMEM2WBReg <= _pipMEM2WBReg_T; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_dataOut_rdata_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      exu_io_dataOut_rdata_r <= io_dataIO_data_read; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      pipWB2ENDWire_r <= 70'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      pipWB2ENDWire_r <= _pipWB2ENDWire_T; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  pipEX2MEMReg = _RAND_0[248:0];
  _RAND_1 = {14{`RANDOM}};
  pipID2ExReg = _RAND_1[430:0];
  _RAND_2 = {1{`RANDOM}};
  pipCSRReg = _RAND_2[8:0];
  _RAND_3 = {5{`RANDOM}};
  pipIF2IDReg = _RAND_3[129:0];
  _RAND_4 = {6{`RANDOM}};
  pipMEM2WBReg = _RAND_4[173:0];
  _RAND_5 = {2{`RANDOM}};
  exu_io_dataOut_rdata_r = _RAND_5[63:0];
  _RAND_6 = {3{`RANDOM}};
  pipWB2ENDWire_r = _RAND_6[69:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Icache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output [31:0]  io_cacheOut_w_addr_o,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [31:0]  io_cacheIn_addr,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          updataICache_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] offset = io_cacheIn_addr[3:0]; // @[Cache.scala 27:31]
  wire [5:0] index = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  wire [21:0] tag = io_cacheIn_addr[31:10]; // @[Cache.scala 29:28]
  reg  cacheState; // @[Cache.scala 32:27]
  wire  _vMuxOut_T_124 = 6'h3f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_63_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_122 = 6'h3e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_62_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_120 = 6'h3d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_61_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_118 = 6'h3c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_60_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_116 = 6'h3b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_59_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_114 = 6'h3a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_58_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_112 = 6'h39 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_57_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_110 = 6'h38 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_56_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_108 = 6'h37 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_55_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_106 = 6'h36 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_54_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_104 = 6'h35 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_53_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_102 = 6'h34 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_52_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_100 = 6'h33 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_51_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_98 = 6'h32 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_50_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_96 = 6'h31 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_49_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_94 = 6'h30 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_48_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_92 = 6'h2f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_47_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_90 = 6'h2e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_46_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_88 = 6'h2d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_45_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_86 = 6'h2c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_44_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_84 = 6'h2b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_43_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_82 = 6'h2a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_42_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_80 = 6'h29 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_41_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_78 = 6'h28 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_40_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_76 = 6'h27 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_39_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_74 = 6'h26 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_38_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_72 = 6'h25 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_37_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_70 = 6'h24 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_36_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_68 = 6'h23 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_35_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_66 = 6'h22 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_34_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_64 = 6'h21 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_33_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_62 = 6'h20 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_32_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_60 = 6'h1f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_31_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_58 = 6'h1e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_30_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_56 = 6'h1d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_29_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_54 = 6'h1c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_28_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_52 = 6'h1b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_27_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_50 = 6'h1a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_26_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_48 = 6'h19 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_25_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_46 = 6'h18 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_24_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_44 = 6'h17 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_23_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_42 = 6'h16 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_22_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_40 = 6'h15 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_21_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_38 = 6'h14 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_20_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_36 = 6'h13 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_19_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_34 = 6'h12 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_18_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_32 = 6'h11 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_17_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_30 = 6'h10 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_16_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_28 = 6'hf == index; // @[Mux.scala 80:60]
  reg  vArrayWire_15_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_26 = 6'he == index; // @[Mux.scala 80:60]
  reg  vArrayWire_14_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_24 = 6'hd == index; // @[Mux.scala 80:60]
  reg  vArrayWire_13_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_22 = 6'hc == index; // @[Mux.scala 80:60]
  reg  vArrayWire_12_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_20 = 6'hb == index; // @[Mux.scala 80:60]
  reg  vArrayWire_11_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_18 = 6'ha == index; // @[Mux.scala 80:60]
  reg  vArrayWire_10_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_16 = 6'h9 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_9_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_14 = 6'h8 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_8_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_12 = 6'h7 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_7_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_10 = 6'h6 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_6_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_8 = 6'h5 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_5_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_6 = 6'h4 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_4_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_4 = 6'h3 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_3_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_2 = 6'h2 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_2_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T = 6'h1 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_1_0_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_0 = 6'h1 == index ? vArrayWire_1_0_r : vArrayWire_0_0_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_0 = 6'h2 == index ? vArrayWire_2_0_r : _vMuxOut_T_1_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_0 = 6'h3 == index ? vArrayWire_3_0_r : _vMuxOut_T_3_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_0 = 6'h4 == index ? vArrayWire_4_0_r : _vMuxOut_T_5_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_0 = 6'h5 == index ? vArrayWire_5_0_r : _vMuxOut_T_7_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_0 = 6'h6 == index ? vArrayWire_6_0_r : _vMuxOut_T_9_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_0 = 6'h7 == index ? vArrayWire_7_0_r : _vMuxOut_T_11_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_0 = 6'h8 == index ? vArrayWire_8_0_r : _vMuxOut_T_13_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_0 = 6'h9 == index ? vArrayWire_9_0_r : _vMuxOut_T_15_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_0 = 6'ha == index ? vArrayWire_10_0_r : _vMuxOut_T_17_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_0 = 6'hb == index ? vArrayWire_11_0_r : _vMuxOut_T_19_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_0 = 6'hc == index ? vArrayWire_12_0_r : _vMuxOut_T_21_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_0 = 6'hd == index ? vArrayWire_13_0_r : _vMuxOut_T_23_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_0 = 6'he == index ? vArrayWire_14_0_r : _vMuxOut_T_25_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_0 = 6'hf == index ? vArrayWire_15_0_r : _vMuxOut_T_27_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_0 = 6'h10 == index ? vArrayWire_16_0_r : _vMuxOut_T_29_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_0 = 6'h11 == index ? vArrayWire_17_0_r : _vMuxOut_T_31_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_0 = 6'h12 == index ? vArrayWire_18_0_r : _vMuxOut_T_33_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_0 = 6'h13 == index ? vArrayWire_19_0_r : _vMuxOut_T_35_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_0 = 6'h14 == index ? vArrayWire_20_0_r : _vMuxOut_T_37_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_0 = 6'h15 == index ? vArrayWire_21_0_r : _vMuxOut_T_39_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_0 = 6'h16 == index ? vArrayWire_22_0_r : _vMuxOut_T_41_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_0 = 6'h17 == index ? vArrayWire_23_0_r : _vMuxOut_T_43_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_0 = 6'h18 == index ? vArrayWire_24_0_r : _vMuxOut_T_45_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_0 = 6'h19 == index ? vArrayWire_25_0_r : _vMuxOut_T_47_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_0 = 6'h1a == index ? vArrayWire_26_0_r : _vMuxOut_T_49_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_0 = 6'h1b == index ? vArrayWire_27_0_r : _vMuxOut_T_51_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_0 = 6'h1c == index ? vArrayWire_28_0_r : _vMuxOut_T_53_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_0 = 6'h1d == index ? vArrayWire_29_0_r : _vMuxOut_T_55_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_0 = 6'h1e == index ? vArrayWire_30_0_r : _vMuxOut_T_57_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_0 = 6'h1f == index ? vArrayWire_31_0_r : _vMuxOut_T_59_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_0 = 6'h20 == index ? vArrayWire_32_0_r : _vMuxOut_T_61_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_0 = 6'h21 == index ? vArrayWire_33_0_r : _vMuxOut_T_63_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_0 = 6'h22 == index ? vArrayWire_34_0_r : _vMuxOut_T_65_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_0 = 6'h23 == index ? vArrayWire_35_0_r : _vMuxOut_T_67_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_0 = 6'h24 == index ? vArrayWire_36_0_r : _vMuxOut_T_69_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_0 = 6'h25 == index ? vArrayWire_37_0_r : _vMuxOut_T_71_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_0 = 6'h26 == index ? vArrayWire_38_0_r : _vMuxOut_T_73_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_0 = 6'h27 == index ? vArrayWire_39_0_r : _vMuxOut_T_75_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_0 = 6'h28 == index ? vArrayWire_40_0_r : _vMuxOut_T_77_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_0 = 6'h29 == index ? vArrayWire_41_0_r : _vMuxOut_T_79_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_0 = 6'h2a == index ? vArrayWire_42_0_r : _vMuxOut_T_81_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_0 = 6'h2b == index ? vArrayWire_43_0_r : _vMuxOut_T_83_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_0 = 6'h2c == index ? vArrayWire_44_0_r : _vMuxOut_T_85_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_0 = 6'h2d == index ? vArrayWire_45_0_r : _vMuxOut_T_87_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_0 = 6'h2e == index ? vArrayWire_46_0_r : _vMuxOut_T_89_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_0 = 6'h2f == index ? vArrayWire_47_0_r : _vMuxOut_T_91_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_0 = 6'h30 == index ? vArrayWire_48_0_r : _vMuxOut_T_93_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_0 = 6'h31 == index ? vArrayWire_49_0_r : _vMuxOut_T_95_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_0 = 6'h32 == index ? vArrayWire_50_0_r : _vMuxOut_T_97_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_0 = 6'h33 == index ? vArrayWire_51_0_r : _vMuxOut_T_99_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_0 = 6'h34 == index ? vArrayWire_52_0_r : _vMuxOut_T_101_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_0 = 6'h35 == index ? vArrayWire_53_0_r : _vMuxOut_T_103_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_0 = 6'h36 == index ? vArrayWire_54_0_r : _vMuxOut_T_105_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_0 = 6'h37 == index ? vArrayWire_55_0_r : _vMuxOut_T_107_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_0 = 6'h38 == index ? vArrayWire_56_0_r : _vMuxOut_T_109_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_0 = 6'h39 == index ? vArrayWire_57_0_r : _vMuxOut_T_111_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_0 = 6'h3a == index ? vArrayWire_58_0_r : _vMuxOut_T_113_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_0 = 6'h3b == index ? vArrayWire_59_0_r : _vMuxOut_T_115_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_0 = 6'h3c == index ? vArrayWire_60_0_r : _vMuxOut_T_117_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_0 = 6'h3d == index ? vArrayWire_61_0_r : _vMuxOut_T_119_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_0 = 6'h3e == index ? vArrayWire_62_0_r : _vMuxOut_T_121_0; // @[Mux.scala 80:57]
  wire  vMuxOut_0 = 6'h3f == index ? vArrayWire_63_0_r : _vMuxOut_T_123_0; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_0_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_0 = 6'h1 == index ? tagArrayWire_1_0_r : tagArrayWire_0_0_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_0 = 6'h2 == index ? tagArrayWire_2_0_r : _tagMuxOut_T_1_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_0 = 6'h3 == index ? tagArrayWire_3_0_r : _tagMuxOut_T_3_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_0 = 6'h4 == index ? tagArrayWire_4_0_r : _tagMuxOut_T_5_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_0 = 6'h5 == index ? tagArrayWire_5_0_r : _tagMuxOut_T_7_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_0 = 6'h6 == index ? tagArrayWire_6_0_r : _tagMuxOut_T_9_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_0 = 6'h7 == index ? tagArrayWire_7_0_r : _tagMuxOut_T_11_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_0 = 6'h8 == index ? tagArrayWire_8_0_r : _tagMuxOut_T_13_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_0 = 6'h9 == index ? tagArrayWire_9_0_r : _tagMuxOut_T_15_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_0 = 6'ha == index ? tagArrayWire_10_0_r : _tagMuxOut_T_17_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_0 = 6'hb == index ? tagArrayWire_11_0_r : _tagMuxOut_T_19_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_0 = 6'hc == index ? tagArrayWire_12_0_r : _tagMuxOut_T_21_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_0 = 6'hd == index ? tagArrayWire_13_0_r : _tagMuxOut_T_23_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_0 = 6'he == index ? tagArrayWire_14_0_r : _tagMuxOut_T_25_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_0 = 6'hf == index ? tagArrayWire_15_0_r : _tagMuxOut_T_27_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_0 = 6'h10 == index ? tagArrayWire_16_0_r : _tagMuxOut_T_29_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_0 = 6'h11 == index ? tagArrayWire_17_0_r : _tagMuxOut_T_31_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_0 = 6'h12 == index ? tagArrayWire_18_0_r : _tagMuxOut_T_33_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_0 = 6'h13 == index ? tagArrayWire_19_0_r : _tagMuxOut_T_35_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_0 = 6'h14 == index ? tagArrayWire_20_0_r : _tagMuxOut_T_37_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_0 = 6'h15 == index ? tagArrayWire_21_0_r : _tagMuxOut_T_39_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_0 = 6'h16 == index ? tagArrayWire_22_0_r : _tagMuxOut_T_41_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_0 = 6'h17 == index ? tagArrayWire_23_0_r : _tagMuxOut_T_43_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_0 = 6'h18 == index ? tagArrayWire_24_0_r : _tagMuxOut_T_45_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_0 = 6'h19 == index ? tagArrayWire_25_0_r : _tagMuxOut_T_47_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_0 = 6'h1a == index ? tagArrayWire_26_0_r : _tagMuxOut_T_49_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_0 = 6'h1b == index ? tagArrayWire_27_0_r : _tagMuxOut_T_51_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_0 = 6'h1c == index ? tagArrayWire_28_0_r : _tagMuxOut_T_53_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_0 = 6'h1d == index ? tagArrayWire_29_0_r : _tagMuxOut_T_55_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_0 = 6'h1e == index ? tagArrayWire_30_0_r : _tagMuxOut_T_57_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_0 = 6'h1f == index ? tagArrayWire_31_0_r : _tagMuxOut_T_59_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_0 = 6'h20 == index ? tagArrayWire_32_0_r : _tagMuxOut_T_61_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_0 = 6'h21 == index ? tagArrayWire_33_0_r : _tagMuxOut_T_63_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_0 = 6'h22 == index ? tagArrayWire_34_0_r : _tagMuxOut_T_65_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_0 = 6'h23 == index ? tagArrayWire_35_0_r : _tagMuxOut_T_67_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_0 = 6'h24 == index ? tagArrayWire_36_0_r : _tagMuxOut_T_69_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_0 = 6'h25 == index ? tagArrayWire_37_0_r : _tagMuxOut_T_71_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_0 = 6'h26 == index ? tagArrayWire_38_0_r : _tagMuxOut_T_73_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_0 = 6'h27 == index ? tagArrayWire_39_0_r : _tagMuxOut_T_75_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_0 = 6'h28 == index ? tagArrayWire_40_0_r : _tagMuxOut_T_77_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_0 = 6'h29 == index ? tagArrayWire_41_0_r : _tagMuxOut_T_79_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_0 = 6'h2a == index ? tagArrayWire_42_0_r : _tagMuxOut_T_81_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_0 = 6'h2b == index ? tagArrayWire_43_0_r : _tagMuxOut_T_83_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_0 = 6'h2c == index ? tagArrayWire_44_0_r : _tagMuxOut_T_85_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_0 = 6'h2d == index ? tagArrayWire_45_0_r : _tagMuxOut_T_87_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_0 = 6'h2e == index ? tagArrayWire_46_0_r : _tagMuxOut_T_89_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_0 = 6'h2f == index ? tagArrayWire_47_0_r : _tagMuxOut_T_91_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_0 = 6'h30 == index ? tagArrayWire_48_0_r : _tagMuxOut_T_93_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_0 = 6'h31 == index ? tagArrayWire_49_0_r : _tagMuxOut_T_95_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_0 = 6'h32 == index ? tagArrayWire_50_0_r : _tagMuxOut_T_97_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_0 = 6'h33 == index ? tagArrayWire_51_0_r : _tagMuxOut_T_99_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_0 = 6'h34 == index ? tagArrayWire_52_0_r : _tagMuxOut_T_101_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_0 = 6'h35 == index ? tagArrayWire_53_0_r : _tagMuxOut_T_103_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_0 = 6'h36 == index ? tagArrayWire_54_0_r : _tagMuxOut_T_105_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_0 = 6'h37 == index ? tagArrayWire_55_0_r : _tagMuxOut_T_107_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_0 = 6'h38 == index ? tagArrayWire_56_0_r : _tagMuxOut_T_109_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_0 = 6'h39 == index ? tagArrayWire_57_0_r : _tagMuxOut_T_111_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_0 = 6'h3a == index ? tagArrayWire_58_0_r : _tagMuxOut_T_113_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_0 = 6'h3b == index ? tagArrayWire_59_0_r : _tagMuxOut_T_115_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_0 = 6'h3c == index ? tagArrayWire_60_0_r : _tagMuxOut_T_117_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_0 = 6'h3d == index ? tagArrayWire_61_0_r : _tagMuxOut_T_119_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_0 = 6'h3e == index ? tagArrayWire_62_0_r : _tagMuxOut_T_121_0; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_0 = 6'h3f == index ? tagArrayWire_63_0_r : _tagMuxOut_T_123_0; // @[Mux.scala 80:57]
  wire  hitArray_0 = vMuxOut_0 & tagMuxOut_0 == tag; // @[Cache.scala 72:60]
  reg  vArrayWire_63_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_1_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_1 = 6'h1 == index ? vArrayWire_1_1_r : vArrayWire_0_1_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_1 = 6'h2 == index ? vArrayWire_2_1_r : _vMuxOut_T_1_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_1 = 6'h3 == index ? vArrayWire_3_1_r : _vMuxOut_T_3_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_1 = 6'h4 == index ? vArrayWire_4_1_r : _vMuxOut_T_5_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_1 = 6'h5 == index ? vArrayWire_5_1_r : _vMuxOut_T_7_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_1 = 6'h6 == index ? vArrayWire_6_1_r : _vMuxOut_T_9_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_1 = 6'h7 == index ? vArrayWire_7_1_r : _vMuxOut_T_11_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_1 = 6'h8 == index ? vArrayWire_8_1_r : _vMuxOut_T_13_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_1 = 6'h9 == index ? vArrayWire_9_1_r : _vMuxOut_T_15_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_1 = 6'ha == index ? vArrayWire_10_1_r : _vMuxOut_T_17_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_1 = 6'hb == index ? vArrayWire_11_1_r : _vMuxOut_T_19_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_1 = 6'hc == index ? vArrayWire_12_1_r : _vMuxOut_T_21_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_1 = 6'hd == index ? vArrayWire_13_1_r : _vMuxOut_T_23_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_1 = 6'he == index ? vArrayWire_14_1_r : _vMuxOut_T_25_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_1 = 6'hf == index ? vArrayWire_15_1_r : _vMuxOut_T_27_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_1 = 6'h10 == index ? vArrayWire_16_1_r : _vMuxOut_T_29_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_1 = 6'h11 == index ? vArrayWire_17_1_r : _vMuxOut_T_31_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_1 = 6'h12 == index ? vArrayWire_18_1_r : _vMuxOut_T_33_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_1 = 6'h13 == index ? vArrayWire_19_1_r : _vMuxOut_T_35_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_1 = 6'h14 == index ? vArrayWire_20_1_r : _vMuxOut_T_37_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_1 = 6'h15 == index ? vArrayWire_21_1_r : _vMuxOut_T_39_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_1 = 6'h16 == index ? vArrayWire_22_1_r : _vMuxOut_T_41_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_1 = 6'h17 == index ? vArrayWire_23_1_r : _vMuxOut_T_43_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_1 = 6'h18 == index ? vArrayWire_24_1_r : _vMuxOut_T_45_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_1 = 6'h19 == index ? vArrayWire_25_1_r : _vMuxOut_T_47_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_1 = 6'h1a == index ? vArrayWire_26_1_r : _vMuxOut_T_49_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_1 = 6'h1b == index ? vArrayWire_27_1_r : _vMuxOut_T_51_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_1 = 6'h1c == index ? vArrayWire_28_1_r : _vMuxOut_T_53_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_1 = 6'h1d == index ? vArrayWire_29_1_r : _vMuxOut_T_55_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_1 = 6'h1e == index ? vArrayWire_30_1_r : _vMuxOut_T_57_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_1 = 6'h1f == index ? vArrayWire_31_1_r : _vMuxOut_T_59_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_1 = 6'h20 == index ? vArrayWire_32_1_r : _vMuxOut_T_61_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_1 = 6'h21 == index ? vArrayWire_33_1_r : _vMuxOut_T_63_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_1 = 6'h22 == index ? vArrayWire_34_1_r : _vMuxOut_T_65_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_1 = 6'h23 == index ? vArrayWire_35_1_r : _vMuxOut_T_67_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_1 = 6'h24 == index ? vArrayWire_36_1_r : _vMuxOut_T_69_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_1 = 6'h25 == index ? vArrayWire_37_1_r : _vMuxOut_T_71_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_1 = 6'h26 == index ? vArrayWire_38_1_r : _vMuxOut_T_73_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_1 = 6'h27 == index ? vArrayWire_39_1_r : _vMuxOut_T_75_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_1 = 6'h28 == index ? vArrayWire_40_1_r : _vMuxOut_T_77_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_1 = 6'h29 == index ? vArrayWire_41_1_r : _vMuxOut_T_79_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_1 = 6'h2a == index ? vArrayWire_42_1_r : _vMuxOut_T_81_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_1 = 6'h2b == index ? vArrayWire_43_1_r : _vMuxOut_T_83_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_1 = 6'h2c == index ? vArrayWire_44_1_r : _vMuxOut_T_85_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_1 = 6'h2d == index ? vArrayWire_45_1_r : _vMuxOut_T_87_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_1 = 6'h2e == index ? vArrayWire_46_1_r : _vMuxOut_T_89_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_1 = 6'h2f == index ? vArrayWire_47_1_r : _vMuxOut_T_91_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_1 = 6'h30 == index ? vArrayWire_48_1_r : _vMuxOut_T_93_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_1 = 6'h31 == index ? vArrayWire_49_1_r : _vMuxOut_T_95_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_1 = 6'h32 == index ? vArrayWire_50_1_r : _vMuxOut_T_97_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_1 = 6'h33 == index ? vArrayWire_51_1_r : _vMuxOut_T_99_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_1 = 6'h34 == index ? vArrayWire_52_1_r : _vMuxOut_T_101_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_1 = 6'h35 == index ? vArrayWire_53_1_r : _vMuxOut_T_103_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_1 = 6'h36 == index ? vArrayWire_54_1_r : _vMuxOut_T_105_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_1 = 6'h37 == index ? vArrayWire_55_1_r : _vMuxOut_T_107_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_1 = 6'h38 == index ? vArrayWire_56_1_r : _vMuxOut_T_109_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_1 = 6'h39 == index ? vArrayWire_57_1_r : _vMuxOut_T_111_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_1 = 6'h3a == index ? vArrayWire_58_1_r : _vMuxOut_T_113_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_1 = 6'h3b == index ? vArrayWire_59_1_r : _vMuxOut_T_115_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_1 = 6'h3c == index ? vArrayWire_60_1_r : _vMuxOut_T_117_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_1 = 6'h3d == index ? vArrayWire_61_1_r : _vMuxOut_T_119_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_1 = 6'h3e == index ? vArrayWire_62_1_r : _vMuxOut_T_121_1; // @[Mux.scala 80:57]
  wire  vMuxOut_1 = 6'h3f == index ? vArrayWire_63_1_r : _vMuxOut_T_123_1; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_1_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_1 = 6'h1 == index ? tagArrayWire_1_1_r : tagArrayWire_0_1_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_1 = 6'h2 == index ? tagArrayWire_2_1_r : _tagMuxOut_T_1_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_1 = 6'h3 == index ? tagArrayWire_3_1_r : _tagMuxOut_T_3_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_1 = 6'h4 == index ? tagArrayWire_4_1_r : _tagMuxOut_T_5_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_1 = 6'h5 == index ? tagArrayWire_5_1_r : _tagMuxOut_T_7_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_1 = 6'h6 == index ? tagArrayWire_6_1_r : _tagMuxOut_T_9_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_1 = 6'h7 == index ? tagArrayWire_7_1_r : _tagMuxOut_T_11_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_1 = 6'h8 == index ? tagArrayWire_8_1_r : _tagMuxOut_T_13_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_1 = 6'h9 == index ? tagArrayWire_9_1_r : _tagMuxOut_T_15_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_1 = 6'ha == index ? tagArrayWire_10_1_r : _tagMuxOut_T_17_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_1 = 6'hb == index ? tagArrayWire_11_1_r : _tagMuxOut_T_19_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_1 = 6'hc == index ? tagArrayWire_12_1_r : _tagMuxOut_T_21_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_1 = 6'hd == index ? tagArrayWire_13_1_r : _tagMuxOut_T_23_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_1 = 6'he == index ? tagArrayWire_14_1_r : _tagMuxOut_T_25_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_1 = 6'hf == index ? tagArrayWire_15_1_r : _tagMuxOut_T_27_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_1 = 6'h10 == index ? tagArrayWire_16_1_r : _tagMuxOut_T_29_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_1 = 6'h11 == index ? tagArrayWire_17_1_r : _tagMuxOut_T_31_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_1 = 6'h12 == index ? tagArrayWire_18_1_r : _tagMuxOut_T_33_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_1 = 6'h13 == index ? tagArrayWire_19_1_r : _tagMuxOut_T_35_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_1 = 6'h14 == index ? tagArrayWire_20_1_r : _tagMuxOut_T_37_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_1 = 6'h15 == index ? tagArrayWire_21_1_r : _tagMuxOut_T_39_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_1 = 6'h16 == index ? tagArrayWire_22_1_r : _tagMuxOut_T_41_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_1 = 6'h17 == index ? tagArrayWire_23_1_r : _tagMuxOut_T_43_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_1 = 6'h18 == index ? tagArrayWire_24_1_r : _tagMuxOut_T_45_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_1 = 6'h19 == index ? tagArrayWire_25_1_r : _tagMuxOut_T_47_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_1 = 6'h1a == index ? tagArrayWire_26_1_r : _tagMuxOut_T_49_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_1 = 6'h1b == index ? tagArrayWire_27_1_r : _tagMuxOut_T_51_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_1 = 6'h1c == index ? tagArrayWire_28_1_r : _tagMuxOut_T_53_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_1 = 6'h1d == index ? tagArrayWire_29_1_r : _tagMuxOut_T_55_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_1 = 6'h1e == index ? tagArrayWire_30_1_r : _tagMuxOut_T_57_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_1 = 6'h1f == index ? tagArrayWire_31_1_r : _tagMuxOut_T_59_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_1 = 6'h20 == index ? tagArrayWire_32_1_r : _tagMuxOut_T_61_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_1 = 6'h21 == index ? tagArrayWire_33_1_r : _tagMuxOut_T_63_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_1 = 6'h22 == index ? tagArrayWire_34_1_r : _tagMuxOut_T_65_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_1 = 6'h23 == index ? tagArrayWire_35_1_r : _tagMuxOut_T_67_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_1 = 6'h24 == index ? tagArrayWire_36_1_r : _tagMuxOut_T_69_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_1 = 6'h25 == index ? tagArrayWire_37_1_r : _tagMuxOut_T_71_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_1 = 6'h26 == index ? tagArrayWire_38_1_r : _tagMuxOut_T_73_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_1 = 6'h27 == index ? tagArrayWire_39_1_r : _tagMuxOut_T_75_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_1 = 6'h28 == index ? tagArrayWire_40_1_r : _tagMuxOut_T_77_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_1 = 6'h29 == index ? tagArrayWire_41_1_r : _tagMuxOut_T_79_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_1 = 6'h2a == index ? tagArrayWire_42_1_r : _tagMuxOut_T_81_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_1 = 6'h2b == index ? tagArrayWire_43_1_r : _tagMuxOut_T_83_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_1 = 6'h2c == index ? tagArrayWire_44_1_r : _tagMuxOut_T_85_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_1 = 6'h2d == index ? tagArrayWire_45_1_r : _tagMuxOut_T_87_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_1 = 6'h2e == index ? tagArrayWire_46_1_r : _tagMuxOut_T_89_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_1 = 6'h2f == index ? tagArrayWire_47_1_r : _tagMuxOut_T_91_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_1 = 6'h30 == index ? tagArrayWire_48_1_r : _tagMuxOut_T_93_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_1 = 6'h31 == index ? tagArrayWire_49_1_r : _tagMuxOut_T_95_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_1 = 6'h32 == index ? tagArrayWire_50_1_r : _tagMuxOut_T_97_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_1 = 6'h33 == index ? tagArrayWire_51_1_r : _tagMuxOut_T_99_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_1 = 6'h34 == index ? tagArrayWire_52_1_r : _tagMuxOut_T_101_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_1 = 6'h35 == index ? tagArrayWire_53_1_r : _tagMuxOut_T_103_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_1 = 6'h36 == index ? tagArrayWire_54_1_r : _tagMuxOut_T_105_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_1 = 6'h37 == index ? tagArrayWire_55_1_r : _tagMuxOut_T_107_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_1 = 6'h38 == index ? tagArrayWire_56_1_r : _tagMuxOut_T_109_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_1 = 6'h39 == index ? tagArrayWire_57_1_r : _tagMuxOut_T_111_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_1 = 6'h3a == index ? tagArrayWire_58_1_r : _tagMuxOut_T_113_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_1 = 6'h3b == index ? tagArrayWire_59_1_r : _tagMuxOut_T_115_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_1 = 6'h3c == index ? tagArrayWire_60_1_r : _tagMuxOut_T_117_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_1 = 6'h3d == index ? tagArrayWire_61_1_r : _tagMuxOut_T_119_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_1 = 6'h3e == index ? tagArrayWire_62_1_r : _tagMuxOut_T_121_1; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_1 = 6'h3f == index ? tagArrayWire_63_1_r : _tagMuxOut_T_123_1; // @[Mux.scala 80:57]
  wire  hitArray_1 = vMuxOut_1 & tagMuxOut_1 == tag; // @[Cache.scala 72:60]
  reg  vArrayWire_63_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_2_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_2 = 6'h1 == index ? vArrayWire_1_2_r : vArrayWire_0_2_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_2 = 6'h2 == index ? vArrayWire_2_2_r : _vMuxOut_T_1_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_2 = 6'h3 == index ? vArrayWire_3_2_r : _vMuxOut_T_3_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_2 = 6'h4 == index ? vArrayWire_4_2_r : _vMuxOut_T_5_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_2 = 6'h5 == index ? vArrayWire_5_2_r : _vMuxOut_T_7_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_2 = 6'h6 == index ? vArrayWire_6_2_r : _vMuxOut_T_9_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_2 = 6'h7 == index ? vArrayWire_7_2_r : _vMuxOut_T_11_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_2 = 6'h8 == index ? vArrayWire_8_2_r : _vMuxOut_T_13_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_2 = 6'h9 == index ? vArrayWire_9_2_r : _vMuxOut_T_15_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_2 = 6'ha == index ? vArrayWire_10_2_r : _vMuxOut_T_17_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_2 = 6'hb == index ? vArrayWire_11_2_r : _vMuxOut_T_19_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_2 = 6'hc == index ? vArrayWire_12_2_r : _vMuxOut_T_21_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_2 = 6'hd == index ? vArrayWire_13_2_r : _vMuxOut_T_23_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_2 = 6'he == index ? vArrayWire_14_2_r : _vMuxOut_T_25_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_2 = 6'hf == index ? vArrayWire_15_2_r : _vMuxOut_T_27_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_2 = 6'h10 == index ? vArrayWire_16_2_r : _vMuxOut_T_29_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_2 = 6'h11 == index ? vArrayWire_17_2_r : _vMuxOut_T_31_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_2 = 6'h12 == index ? vArrayWire_18_2_r : _vMuxOut_T_33_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_2 = 6'h13 == index ? vArrayWire_19_2_r : _vMuxOut_T_35_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_2 = 6'h14 == index ? vArrayWire_20_2_r : _vMuxOut_T_37_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_2 = 6'h15 == index ? vArrayWire_21_2_r : _vMuxOut_T_39_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_2 = 6'h16 == index ? vArrayWire_22_2_r : _vMuxOut_T_41_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_2 = 6'h17 == index ? vArrayWire_23_2_r : _vMuxOut_T_43_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_2 = 6'h18 == index ? vArrayWire_24_2_r : _vMuxOut_T_45_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_2 = 6'h19 == index ? vArrayWire_25_2_r : _vMuxOut_T_47_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_2 = 6'h1a == index ? vArrayWire_26_2_r : _vMuxOut_T_49_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_2 = 6'h1b == index ? vArrayWire_27_2_r : _vMuxOut_T_51_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_2 = 6'h1c == index ? vArrayWire_28_2_r : _vMuxOut_T_53_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_2 = 6'h1d == index ? vArrayWire_29_2_r : _vMuxOut_T_55_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_2 = 6'h1e == index ? vArrayWire_30_2_r : _vMuxOut_T_57_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_2 = 6'h1f == index ? vArrayWire_31_2_r : _vMuxOut_T_59_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_2 = 6'h20 == index ? vArrayWire_32_2_r : _vMuxOut_T_61_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_2 = 6'h21 == index ? vArrayWire_33_2_r : _vMuxOut_T_63_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_2 = 6'h22 == index ? vArrayWire_34_2_r : _vMuxOut_T_65_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_2 = 6'h23 == index ? vArrayWire_35_2_r : _vMuxOut_T_67_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_2 = 6'h24 == index ? vArrayWire_36_2_r : _vMuxOut_T_69_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_2 = 6'h25 == index ? vArrayWire_37_2_r : _vMuxOut_T_71_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_2 = 6'h26 == index ? vArrayWire_38_2_r : _vMuxOut_T_73_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_2 = 6'h27 == index ? vArrayWire_39_2_r : _vMuxOut_T_75_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_2 = 6'h28 == index ? vArrayWire_40_2_r : _vMuxOut_T_77_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_2 = 6'h29 == index ? vArrayWire_41_2_r : _vMuxOut_T_79_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_2 = 6'h2a == index ? vArrayWire_42_2_r : _vMuxOut_T_81_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_2 = 6'h2b == index ? vArrayWire_43_2_r : _vMuxOut_T_83_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_2 = 6'h2c == index ? vArrayWire_44_2_r : _vMuxOut_T_85_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_2 = 6'h2d == index ? vArrayWire_45_2_r : _vMuxOut_T_87_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_2 = 6'h2e == index ? vArrayWire_46_2_r : _vMuxOut_T_89_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_2 = 6'h2f == index ? vArrayWire_47_2_r : _vMuxOut_T_91_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_2 = 6'h30 == index ? vArrayWire_48_2_r : _vMuxOut_T_93_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_2 = 6'h31 == index ? vArrayWire_49_2_r : _vMuxOut_T_95_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_2 = 6'h32 == index ? vArrayWire_50_2_r : _vMuxOut_T_97_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_2 = 6'h33 == index ? vArrayWire_51_2_r : _vMuxOut_T_99_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_2 = 6'h34 == index ? vArrayWire_52_2_r : _vMuxOut_T_101_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_2 = 6'h35 == index ? vArrayWire_53_2_r : _vMuxOut_T_103_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_2 = 6'h36 == index ? vArrayWire_54_2_r : _vMuxOut_T_105_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_2 = 6'h37 == index ? vArrayWire_55_2_r : _vMuxOut_T_107_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_2 = 6'h38 == index ? vArrayWire_56_2_r : _vMuxOut_T_109_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_2 = 6'h39 == index ? vArrayWire_57_2_r : _vMuxOut_T_111_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_2 = 6'h3a == index ? vArrayWire_58_2_r : _vMuxOut_T_113_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_2 = 6'h3b == index ? vArrayWire_59_2_r : _vMuxOut_T_115_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_2 = 6'h3c == index ? vArrayWire_60_2_r : _vMuxOut_T_117_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_2 = 6'h3d == index ? vArrayWire_61_2_r : _vMuxOut_T_119_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_2 = 6'h3e == index ? vArrayWire_62_2_r : _vMuxOut_T_121_2; // @[Mux.scala 80:57]
  wire  vMuxOut_2 = 6'h3f == index ? vArrayWire_63_2_r : _vMuxOut_T_123_2; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_2_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_2 = 6'h1 == index ? tagArrayWire_1_2_r : tagArrayWire_0_2_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_2 = 6'h2 == index ? tagArrayWire_2_2_r : _tagMuxOut_T_1_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_2 = 6'h3 == index ? tagArrayWire_3_2_r : _tagMuxOut_T_3_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_2 = 6'h4 == index ? tagArrayWire_4_2_r : _tagMuxOut_T_5_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_2 = 6'h5 == index ? tagArrayWire_5_2_r : _tagMuxOut_T_7_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_2 = 6'h6 == index ? tagArrayWire_6_2_r : _tagMuxOut_T_9_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_2 = 6'h7 == index ? tagArrayWire_7_2_r : _tagMuxOut_T_11_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_2 = 6'h8 == index ? tagArrayWire_8_2_r : _tagMuxOut_T_13_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_2 = 6'h9 == index ? tagArrayWire_9_2_r : _tagMuxOut_T_15_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_2 = 6'ha == index ? tagArrayWire_10_2_r : _tagMuxOut_T_17_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_2 = 6'hb == index ? tagArrayWire_11_2_r : _tagMuxOut_T_19_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_2 = 6'hc == index ? tagArrayWire_12_2_r : _tagMuxOut_T_21_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_2 = 6'hd == index ? tagArrayWire_13_2_r : _tagMuxOut_T_23_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_2 = 6'he == index ? tagArrayWire_14_2_r : _tagMuxOut_T_25_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_2 = 6'hf == index ? tagArrayWire_15_2_r : _tagMuxOut_T_27_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_2 = 6'h10 == index ? tagArrayWire_16_2_r : _tagMuxOut_T_29_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_2 = 6'h11 == index ? tagArrayWire_17_2_r : _tagMuxOut_T_31_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_2 = 6'h12 == index ? tagArrayWire_18_2_r : _tagMuxOut_T_33_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_2 = 6'h13 == index ? tagArrayWire_19_2_r : _tagMuxOut_T_35_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_2 = 6'h14 == index ? tagArrayWire_20_2_r : _tagMuxOut_T_37_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_2 = 6'h15 == index ? tagArrayWire_21_2_r : _tagMuxOut_T_39_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_2 = 6'h16 == index ? tagArrayWire_22_2_r : _tagMuxOut_T_41_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_2 = 6'h17 == index ? tagArrayWire_23_2_r : _tagMuxOut_T_43_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_2 = 6'h18 == index ? tagArrayWire_24_2_r : _tagMuxOut_T_45_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_2 = 6'h19 == index ? tagArrayWire_25_2_r : _tagMuxOut_T_47_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_2 = 6'h1a == index ? tagArrayWire_26_2_r : _tagMuxOut_T_49_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_2 = 6'h1b == index ? tagArrayWire_27_2_r : _tagMuxOut_T_51_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_2 = 6'h1c == index ? tagArrayWire_28_2_r : _tagMuxOut_T_53_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_2 = 6'h1d == index ? tagArrayWire_29_2_r : _tagMuxOut_T_55_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_2 = 6'h1e == index ? tagArrayWire_30_2_r : _tagMuxOut_T_57_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_2 = 6'h1f == index ? tagArrayWire_31_2_r : _tagMuxOut_T_59_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_2 = 6'h20 == index ? tagArrayWire_32_2_r : _tagMuxOut_T_61_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_2 = 6'h21 == index ? tagArrayWire_33_2_r : _tagMuxOut_T_63_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_2 = 6'h22 == index ? tagArrayWire_34_2_r : _tagMuxOut_T_65_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_2 = 6'h23 == index ? tagArrayWire_35_2_r : _tagMuxOut_T_67_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_2 = 6'h24 == index ? tagArrayWire_36_2_r : _tagMuxOut_T_69_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_2 = 6'h25 == index ? tagArrayWire_37_2_r : _tagMuxOut_T_71_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_2 = 6'h26 == index ? tagArrayWire_38_2_r : _tagMuxOut_T_73_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_2 = 6'h27 == index ? tagArrayWire_39_2_r : _tagMuxOut_T_75_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_2 = 6'h28 == index ? tagArrayWire_40_2_r : _tagMuxOut_T_77_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_2 = 6'h29 == index ? tagArrayWire_41_2_r : _tagMuxOut_T_79_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_2 = 6'h2a == index ? tagArrayWire_42_2_r : _tagMuxOut_T_81_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_2 = 6'h2b == index ? tagArrayWire_43_2_r : _tagMuxOut_T_83_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_2 = 6'h2c == index ? tagArrayWire_44_2_r : _tagMuxOut_T_85_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_2 = 6'h2d == index ? tagArrayWire_45_2_r : _tagMuxOut_T_87_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_2 = 6'h2e == index ? tagArrayWire_46_2_r : _tagMuxOut_T_89_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_2 = 6'h2f == index ? tagArrayWire_47_2_r : _tagMuxOut_T_91_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_2 = 6'h30 == index ? tagArrayWire_48_2_r : _tagMuxOut_T_93_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_2 = 6'h31 == index ? tagArrayWire_49_2_r : _tagMuxOut_T_95_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_2 = 6'h32 == index ? tagArrayWire_50_2_r : _tagMuxOut_T_97_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_2 = 6'h33 == index ? tagArrayWire_51_2_r : _tagMuxOut_T_99_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_2 = 6'h34 == index ? tagArrayWire_52_2_r : _tagMuxOut_T_101_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_2 = 6'h35 == index ? tagArrayWire_53_2_r : _tagMuxOut_T_103_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_2 = 6'h36 == index ? tagArrayWire_54_2_r : _tagMuxOut_T_105_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_2 = 6'h37 == index ? tagArrayWire_55_2_r : _tagMuxOut_T_107_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_2 = 6'h38 == index ? tagArrayWire_56_2_r : _tagMuxOut_T_109_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_2 = 6'h39 == index ? tagArrayWire_57_2_r : _tagMuxOut_T_111_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_2 = 6'h3a == index ? tagArrayWire_58_2_r : _tagMuxOut_T_113_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_2 = 6'h3b == index ? tagArrayWire_59_2_r : _tagMuxOut_T_115_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_2 = 6'h3c == index ? tagArrayWire_60_2_r : _tagMuxOut_T_117_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_2 = 6'h3d == index ? tagArrayWire_61_2_r : _tagMuxOut_T_119_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_2 = 6'h3e == index ? tagArrayWire_62_2_r : _tagMuxOut_T_121_2; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_2 = 6'h3f == index ? tagArrayWire_63_2_r : _tagMuxOut_T_123_2; // @[Mux.scala 80:57]
  wire  hitArray_2 = vMuxOut_2 & tagMuxOut_2 == tag; // @[Cache.scala 72:60]
  reg  vArrayWire_63_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_3_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_3 = 6'h1 == index ? vArrayWire_1_3_r : vArrayWire_0_3_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_3 = 6'h2 == index ? vArrayWire_2_3_r : _vMuxOut_T_1_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_3 = 6'h3 == index ? vArrayWire_3_3_r : _vMuxOut_T_3_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_3 = 6'h4 == index ? vArrayWire_4_3_r : _vMuxOut_T_5_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_3 = 6'h5 == index ? vArrayWire_5_3_r : _vMuxOut_T_7_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_3 = 6'h6 == index ? vArrayWire_6_3_r : _vMuxOut_T_9_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_3 = 6'h7 == index ? vArrayWire_7_3_r : _vMuxOut_T_11_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_3 = 6'h8 == index ? vArrayWire_8_3_r : _vMuxOut_T_13_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_3 = 6'h9 == index ? vArrayWire_9_3_r : _vMuxOut_T_15_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_3 = 6'ha == index ? vArrayWire_10_3_r : _vMuxOut_T_17_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_3 = 6'hb == index ? vArrayWire_11_3_r : _vMuxOut_T_19_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_3 = 6'hc == index ? vArrayWire_12_3_r : _vMuxOut_T_21_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_3 = 6'hd == index ? vArrayWire_13_3_r : _vMuxOut_T_23_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_3 = 6'he == index ? vArrayWire_14_3_r : _vMuxOut_T_25_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_3 = 6'hf == index ? vArrayWire_15_3_r : _vMuxOut_T_27_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_3 = 6'h10 == index ? vArrayWire_16_3_r : _vMuxOut_T_29_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_3 = 6'h11 == index ? vArrayWire_17_3_r : _vMuxOut_T_31_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_3 = 6'h12 == index ? vArrayWire_18_3_r : _vMuxOut_T_33_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_3 = 6'h13 == index ? vArrayWire_19_3_r : _vMuxOut_T_35_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_3 = 6'h14 == index ? vArrayWire_20_3_r : _vMuxOut_T_37_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_3 = 6'h15 == index ? vArrayWire_21_3_r : _vMuxOut_T_39_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_3 = 6'h16 == index ? vArrayWire_22_3_r : _vMuxOut_T_41_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_3 = 6'h17 == index ? vArrayWire_23_3_r : _vMuxOut_T_43_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_3 = 6'h18 == index ? vArrayWire_24_3_r : _vMuxOut_T_45_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_3 = 6'h19 == index ? vArrayWire_25_3_r : _vMuxOut_T_47_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_3 = 6'h1a == index ? vArrayWire_26_3_r : _vMuxOut_T_49_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_3 = 6'h1b == index ? vArrayWire_27_3_r : _vMuxOut_T_51_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_3 = 6'h1c == index ? vArrayWire_28_3_r : _vMuxOut_T_53_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_3 = 6'h1d == index ? vArrayWire_29_3_r : _vMuxOut_T_55_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_3 = 6'h1e == index ? vArrayWire_30_3_r : _vMuxOut_T_57_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_3 = 6'h1f == index ? vArrayWire_31_3_r : _vMuxOut_T_59_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_3 = 6'h20 == index ? vArrayWire_32_3_r : _vMuxOut_T_61_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_3 = 6'h21 == index ? vArrayWire_33_3_r : _vMuxOut_T_63_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_3 = 6'h22 == index ? vArrayWire_34_3_r : _vMuxOut_T_65_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_3 = 6'h23 == index ? vArrayWire_35_3_r : _vMuxOut_T_67_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_3 = 6'h24 == index ? vArrayWire_36_3_r : _vMuxOut_T_69_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_3 = 6'h25 == index ? vArrayWire_37_3_r : _vMuxOut_T_71_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_3 = 6'h26 == index ? vArrayWire_38_3_r : _vMuxOut_T_73_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_3 = 6'h27 == index ? vArrayWire_39_3_r : _vMuxOut_T_75_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_3 = 6'h28 == index ? vArrayWire_40_3_r : _vMuxOut_T_77_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_3 = 6'h29 == index ? vArrayWire_41_3_r : _vMuxOut_T_79_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_3 = 6'h2a == index ? vArrayWire_42_3_r : _vMuxOut_T_81_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_3 = 6'h2b == index ? vArrayWire_43_3_r : _vMuxOut_T_83_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_3 = 6'h2c == index ? vArrayWire_44_3_r : _vMuxOut_T_85_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_3 = 6'h2d == index ? vArrayWire_45_3_r : _vMuxOut_T_87_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_3 = 6'h2e == index ? vArrayWire_46_3_r : _vMuxOut_T_89_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_3 = 6'h2f == index ? vArrayWire_47_3_r : _vMuxOut_T_91_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_3 = 6'h30 == index ? vArrayWire_48_3_r : _vMuxOut_T_93_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_3 = 6'h31 == index ? vArrayWire_49_3_r : _vMuxOut_T_95_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_3 = 6'h32 == index ? vArrayWire_50_3_r : _vMuxOut_T_97_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_3 = 6'h33 == index ? vArrayWire_51_3_r : _vMuxOut_T_99_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_3 = 6'h34 == index ? vArrayWire_52_3_r : _vMuxOut_T_101_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_3 = 6'h35 == index ? vArrayWire_53_3_r : _vMuxOut_T_103_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_3 = 6'h36 == index ? vArrayWire_54_3_r : _vMuxOut_T_105_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_3 = 6'h37 == index ? vArrayWire_55_3_r : _vMuxOut_T_107_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_3 = 6'h38 == index ? vArrayWire_56_3_r : _vMuxOut_T_109_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_3 = 6'h39 == index ? vArrayWire_57_3_r : _vMuxOut_T_111_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_3 = 6'h3a == index ? vArrayWire_58_3_r : _vMuxOut_T_113_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_3 = 6'h3b == index ? vArrayWire_59_3_r : _vMuxOut_T_115_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_3 = 6'h3c == index ? vArrayWire_60_3_r : _vMuxOut_T_117_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_3 = 6'h3d == index ? vArrayWire_61_3_r : _vMuxOut_T_119_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_3 = 6'h3e == index ? vArrayWire_62_3_r : _vMuxOut_T_121_3; // @[Mux.scala 80:57]
  wire  vMuxOut_3 = 6'h3f == index ? vArrayWire_63_3_r : _vMuxOut_T_123_3; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_3_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_3 = 6'h1 == index ? tagArrayWire_1_3_r : tagArrayWire_0_3_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_3 = 6'h2 == index ? tagArrayWire_2_3_r : _tagMuxOut_T_1_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_3 = 6'h3 == index ? tagArrayWire_3_3_r : _tagMuxOut_T_3_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_3 = 6'h4 == index ? tagArrayWire_4_3_r : _tagMuxOut_T_5_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_3 = 6'h5 == index ? tagArrayWire_5_3_r : _tagMuxOut_T_7_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_3 = 6'h6 == index ? tagArrayWire_6_3_r : _tagMuxOut_T_9_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_3 = 6'h7 == index ? tagArrayWire_7_3_r : _tagMuxOut_T_11_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_3 = 6'h8 == index ? tagArrayWire_8_3_r : _tagMuxOut_T_13_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_3 = 6'h9 == index ? tagArrayWire_9_3_r : _tagMuxOut_T_15_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_3 = 6'ha == index ? tagArrayWire_10_3_r : _tagMuxOut_T_17_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_3 = 6'hb == index ? tagArrayWire_11_3_r : _tagMuxOut_T_19_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_3 = 6'hc == index ? tagArrayWire_12_3_r : _tagMuxOut_T_21_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_3 = 6'hd == index ? tagArrayWire_13_3_r : _tagMuxOut_T_23_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_3 = 6'he == index ? tagArrayWire_14_3_r : _tagMuxOut_T_25_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_3 = 6'hf == index ? tagArrayWire_15_3_r : _tagMuxOut_T_27_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_3 = 6'h10 == index ? tagArrayWire_16_3_r : _tagMuxOut_T_29_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_3 = 6'h11 == index ? tagArrayWire_17_3_r : _tagMuxOut_T_31_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_3 = 6'h12 == index ? tagArrayWire_18_3_r : _tagMuxOut_T_33_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_3 = 6'h13 == index ? tagArrayWire_19_3_r : _tagMuxOut_T_35_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_3 = 6'h14 == index ? tagArrayWire_20_3_r : _tagMuxOut_T_37_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_3 = 6'h15 == index ? tagArrayWire_21_3_r : _tagMuxOut_T_39_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_3 = 6'h16 == index ? tagArrayWire_22_3_r : _tagMuxOut_T_41_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_3 = 6'h17 == index ? tagArrayWire_23_3_r : _tagMuxOut_T_43_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_3 = 6'h18 == index ? tagArrayWire_24_3_r : _tagMuxOut_T_45_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_3 = 6'h19 == index ? tagArrayWire_25_3_r : _tagMuxOut_T_47_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_3 = 6'h1a == index ? tagArrayWire_26_3_r : _tagMuxOut_T_49_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_3 = 6'h1b == index ? tagArrayWire_27_3_r : _tagMuxOut_T_51_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_3 = 6'h1c == index ? tagArrayWire_28_3_r : _tagMuxOut_T_53_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_3 = 6'h1d == index ? tagArrayWire_29_3_r : _tagMuxOut_T_55_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_3 = 6'h1e == index ? tagArrayWire_30_3_r : _tagMuxOut_T_57_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_3 = 6'h1f == index ? tagArrayWire_31_3_r : _tagMuxOut_T_59_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_3 = 6'h20 == index ? tagArrayWire_32_3_r : _tagMuxOut_T_61_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_3 = 6'h21 == index ? tagArrayWire_33_3_r : _tagMuxOut_T_63_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_3 = 6'h22 == index ? tagArrayWire_34_3_r : _tagMuxOut_T_65_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_3 = 6'h23 == index ? tagArrayWire_35_3_r : _tagMuxOut_T_67_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_3 = 6'h24 == index ? tagArrayWire_36_3_r : _tagMuxOut_T_69_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_3 = 6'h25 == index ? tagArrayWire_37_3_r : _tagMuxOut_T_71_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_3 = 6'h26 == index ? tagArrayWire_38_3_r : _tagMuxOut_T_73_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_3 = 6'h27 == index ? tagArrayWire_39_3_r : _tagMuxOut_T_75_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_3 = 6'h28 == index ? tagArrayWire_40_3_r : _tagMuxOut_T_77_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_3 = 6'h29 == index ? tagArrayWire_41_3_r : _tagMuxOut_T_79_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_3 = 6'h2a == index ? tagArrayWire_42_3_r : _tagMuxOut_T_81_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_3 = 6'h2b == index ? tagArrayWire_43_3_r : _tagMuxOut_T_83_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_3 = 6'h2c == index ? tagArrayWire_44_3_r : _tagMuxOut_T_85_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_3 = 6'h2d == index ? tagArrayWire_45_3_r : _tagMuxOut_T_87_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_3 = 6'h2e == index ? tagArrayWire_46_3_r : _tagMuxOut_T_89_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_3 = 6'h2f == index ? tagArrayWire_47_3_r : _tagMuxOut_T_91_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_3 = 6'h30 == index ? tagArrayWire_48_3_r : _tagMuxOut_T_93_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_3 = 6'h31 == index ? tagArrayWire_49_3_r : _tagMuxOut_T_95_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_3 = 6'h32 == index ? tagArrayWire_50_3_r : _tagMuxOut_T_97_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_3 = 6'h33 == index ? tagArrayWire_51_3_r : _tagMuxOut_T_99_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_3 = 6'h34 == index ? tagArrayWire_52_3_r : _tagMuxOut_T_101_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_3 = 6'h35 == index ? tagArrayWire_53_3_r : _tagMuxOut_T_103_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_3 = 6'h36 == index ? tagArrayWire_54_3_r : _tagMuxOut_T_105_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_3 = 6'h37 == index ? tagArrayWire_55_3_r : _tagMuxOut_T_107_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_3 = 6'h38 == index ? tagArrayWire_56_3_r : _tagMuxOut_T_109_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_3 = 6'h39 == index ? tagArrayWire_57_3_r : _tagMuxOut_T_111_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_3 = 6'h3a == index ? tagArrayWire_58_3_r : _tagMuxOut_T_113_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_3 = 6'h3b == index ? tagArrayWire_59_3_r : _tagMuxOut_T_115_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_3 = 6'h3c == index ? tagArrayWire_60_3_r : _tagMuxOut_T_117_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_3 = 6'h3d == index ? tagArrayWire_61_3_r : _tagMuxOut_T_119_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_3 = 6'h3e == index ? tagArrayWire_62_3_r : _tagMuxOut_T_121_3; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_3 = 6'h3f == index ? tagArrayWire_63_3_r : _tagMuxOut_T_123_3; // @[Mux.scala 80:57]
  wire  hitArray_3 = vMuxOut_3 & tagMuxOut_3 == tag; // @[Cache.scala 72:60]
  wire  hit = hitArray_0 | hitArray_1 | hitArray_2 | hitArray_3; // @[Cache.scala 73:49]
  wire  IdleMux = io_cacheIn_valid & ~hit; // @[Cache.scala 35:38]
  wire  isIdle = ~cacheState; // @[Cache.scala 45:27]
  wire [127:0] _waysel_T = hitArray_0 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_1 = hitArray_1 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_2 = hitArray_2 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_3 = hitArray_3 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_4 = _waysel_T | _waysel_T_1; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_5 = _waysel_T_4 | _waysel_T_2; // @[Mux.scala 27:72]
  wire [127:0] waysel = _waysel_T_5 | _waysel_T_3; // @[Mux.scala 27:72]
  reg [1:0] selArrayWire_1_r; // @[Reg.scala 27:20]
  reg [1:0] selArrayWire_0_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_1 = 6'h1 == index ? selArrayWire_1_r : selArrayWire_0_r; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_2_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_3 = 6'h2 == index ? selArrayWire_2_r : _sramSel_T_1; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_3_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_5 = 6'h3 == index ? selArrayWire_3_r : _sramSel_T_3; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_4_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_7 = 6'h4 == index ? selArrayWire_4_r : _sramSel_T_5; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_5_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_9 = 6'h5 == index ? selArrayWire_5_r : _sramSel_T_7; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_6_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_11 = 6'h6 == index ? selArrayWire_6_r : _sramSel_T_9; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_7_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_13 = 6'h7 == index ? selArrayWire_7_r : _sramSel_T_11; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_8_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_15 = 6'h8 == index ? selArrayWire_8_r : _sramSel_T_13; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_9_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_17 = 6'h9 == index ? selArrayWire_9_r : _sramSel_T_15; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_10_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_19 = 6'ha == index ? selArrayWire_10_r : _sramSel_T_17; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_11_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_21 = 6'hb == index ? selArrayWire_11_r : _sramSel_T_19; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_12_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_23 = 6'hc == index ? selArrayWire_12_r : _sramSel_T_21; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_13_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_25 = 6'hd == index ? selArrayWire_13_r : _sramSel_T_23; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_14_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_27 = 6'he == index ? selArrayWire_14_r : _sramSel_T_25; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_15_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_29 = 6'hf == index ? selArrayWire_15_r : _sramSel_T_27; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_16_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_31 = 6'h10 == index ? selArrayWire_16_r : _sramSel_T_29; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_17_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_33 = 6'h11 == index ? selArrayWire_17_r : _sramSel_T_31; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_18_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_35 = 6'h12 == index ? selArrayWire_18_r : _sramSel_T_33; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_19_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_37 = 6'h13 == index ? selArrayWire_19_r : _sramSel_T_35; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_20_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_39 = 6'h14 == index ? selArrayWire_20_r : _sramSel_T_37; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_21_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_41 = 6'h15 == index ? selArrayWire_21_r : _sramSel_T_39; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_22_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_43 = 6'h16 == index ? selArrayWire_22_r : _sramSel_T_41; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_23_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_45 = 6'h17 == index ? selArrayWire_23_r : _sramSel_T_43; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_24_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_47 = 6'h18 == index ? selArrayWire_24_r : _sramSel_T_45; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_25_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_49 = 6'h19 == index ? selArrayWire_25_r : _sramSel_T_47; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_26_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_51 = 6'h1a == index ? selArrayWire_26_r : _sramSel_T_49; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_27_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_53 = 6'h1b == index ? selArrayWire_27_r : _sramSel_T_51; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_28_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_55 = 6'h1c == index ? selArrayWire_28_r : _sramSel_T_53; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_29_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_57 = 6'h1d == index ? selArrayWire_29_r : _sramSel_T_55; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_30_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_59 = 6'h1e == index ? selArrayWire_30_r : _sramSel_T_57; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_31_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_61 = 6'h1f == index ? selArrayWire_31_r : _sramSel_T_59; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_32_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_63 = 6'h20 == index ? selArrayWire_32_r : _sramSel_T_61; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_33_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_65 = 6'h21 == index ? selArrayWire_33_r : _sramSel_T_63; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_34_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_67 = 6'h22 == index ? selArrayWire_34_r : _sramSel_T_65; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_35_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_69 = 6'h23 == index ? selArrayWire_35_r : _sramSel_T_67; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_36_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_71 = 6'h24 == index ? selArrayWire_36_r : _sramSel_T_69; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_37_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_73 = 6'h25 == index ? selArrayWire_37_r : _sramSel_T_71; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_38_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_75 = 6'h26 == index ? selArrayWire_38_r : _sramSel_T_73; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_39_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_77 = 6'h27 == index ? selArrayWire_39_r : _sramSel_T_75; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_40_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_79 = 6'h28 == index ? selArrayWire_40_r : _sramSel_T_77; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_41_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_81 = 6'h29 == index ? selArrayWire_41_r : _sramSel_T_79; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_42_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_83 = 6'h2a == index ? selArrayWire_42_r : _sramSel_T_81; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_43_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_85 = 6'h2b == index ? selArrayWire_43_r : _sramSel_T_83; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_44_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_87 = 6'h2c == index ? selArrayWire_44_r : _sramSel_T_85; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_45_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_89 = 6'h2d == index ? selArrayWire_45_r : _sramSel_T_87; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_46_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_91 = 6'h2e == index ? selArrayWire_46_r : _sramSel_T_89; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_47_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_93 = 6'h2f == index ? selArrayWire_47_r : _sramSel_T_91; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_48_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_95 = 6'h30 == index ? selArrayWire_48_r : _sramSel_T_93; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_49_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_97 = 6'h31 == index ? selArrayWire_49_r : _sramSel_T_95; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_50_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_99 = 6'h32 == index ? selArrayWire_50_r : _sramSel_T_97; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_51_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_101 = 6'h33 == index ? selArrayWire_51_r : _sramSel_T_99; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_52_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_103 = 6'h34 == index ? selArrayWire_52_r : _sramSel_T_101; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_53_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_105 = 6'h35 == index ? selArrayWire_53_r : _sramSel_T_103; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_54_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_107 = 6'h36 == index ? selArrayWire_54_r : _sramSel_T_105; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_55_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_109 = 6'h37 == index ? selArrayWire_55_r : _sramSel_T_107; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_56_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_111 = 6'h38 == index ? selArrayWire_56_r : _sramSel_T_109; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_57_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_113 = 6'h39 == index ? selArrayWire_57_r : _sramSel_T_111; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_58_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_115 = 6'h3a == index ? selArrayWire_58_r : _sramSel_T_113; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_59_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_117 = 6'h3b == index ? selArrayWire_59_r : _sramSel_T_115; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_60_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_119 = 6'h3c == index ? selArrayWire_60_r : _sramSel_T_117; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_61_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_121 = 6'h3d == index ? selArrayWire_61_r : _sramSel_T_119; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_62_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_123 = 6'h3e == index ? selArrayWire_62_r : _sramSel_T_121; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_63_r; // @[Reg.scala 27:20]
  wire [1:0] sramSel = 6'h3f == index ? selArrayWire_63_r : _sramSel_T_123; // @[Mux.scala 80:57]
  wire [27:0] io_cacheOut_ar_addr_o_hi = io_cacheIn_addr[31:4]; // @[Cache.scala 104:48]
  wire [1:0] _selArrayWire_0_T_1 = selArrayWire_0_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_0_T_3 = io_cacheOut_r_last_i & 6'h0 == index; // @[Cache.scala 111:28]
  wire  _tagArrayWire_0_0_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _T_1 = reset | updataICache_0; // @[Cache.scala 115:33]
  wire  _GEN_2 = _tagArrayWire_0_0_T_4 | vArrayWire_0_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_1_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_4 = _tagArrayWire_0_1_T_4 | vArrayWire_0_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_2_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_6 = _tagArrayWire_0_2_T_4 | vArrayWire_0_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_3_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_8 = _tagArrayWire_0_3_T_4 | vArrayWire_0_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_1_T_1 = selArrayWire_1_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_1_T_3 = io_cacheOut_r_last_i & _vMuxOut_T; // @[Cache.scala 111:28]
  wire  _tagArrayWire_1_0_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_11 = _tagArrayWire_1_0_T_4 | vArrayWire_1_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_1_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_13 = _tagArrayWire_1_1_T_4 | vArrayWire_1_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_2_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_15 = _tagArrayWire_1_2_T_4 | vArrayWire_1_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_3_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_17 = _tagArrayWire_1_3_T_4 | vArrayWire_1_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_2_T_1 = selArrayWire_2_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_2_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_2; // @[Cache.scala 111:28]
  wire  _tagArrayWire_2_0_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_20 = _tagArrayWire_2_0_T_4 | vArrayWire_2_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_1_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_22 = _tagArrayWire_2_1_T_4 | vArrayWire_2_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_2_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_24 = _tagArrayWire_2_2_T_4 | vArrayWire_2_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_3_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_26 = _tagArrayWire_2_3_T_4 | vArrayWire_2_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_3_T_1 = selArrayWire_3_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_3_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_4; // @[Cache.scala 111:28]
  wire  _tagArrayWire_3_0_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_29 = _tagArrayWire_3_0_T_4 | vArrayWire_3_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_1_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_31 = _tagArrayWire_3_1_T_4 | vArrayWire_3_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_2_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_33 = _tagArrayWire_3_2_T_4 | vArrayWire_3_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_3_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_35 = _tagArrayWire_3_3_T_4 | vArrayWire_3_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_4_T_1 = selArrayWire_4_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_4_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_6; // @[Cache.scala 111:28]
  wire  _tagArrayWire_4_0_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_38 = _tagArrayWire_4_0_T_4 | vArrayWire_4_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_1_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_40 = _tagArrayWire_4_1_T_4 | vArrayWire_4_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_2_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_42 = _tagArrayWire_4_2_T_4 | vArrayWire_4_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_3_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_44 = _tagArrayWire_4_3_T_4 | vArrayWire_4_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_5_T_1 = selArrayWire_5_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_5_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_8; // @[Cache.scala 111:28]
  wire  _tagArrayWire_5_0_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_47 = _tagArrayWire_5_0_T_4 | vArrayWire_5_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_1_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_49 = _tagArrayWire_5_1_T_4 | vArrayWire_5_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_2_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_51 = _tagArrayWire_5_2_T_4 | vArrayWire_5_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_3_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_53 = _tagArrayWire_5_3_T_4 | vArrayWire_5_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_6_T_1 = selArrayWire_6_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_6_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_10; // @[Cache.scala 111:28]
  wire  _tagArrayWire_6_0_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_56 = _tagArrayWire_6_0_T_4 | vArrayWire_6_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_1_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_58 = _tagArrayWire_6_1_T_4 | vArrayWire_6_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_2_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_60 = _tagArrayWire_6_2_T_4 | vArrayWire_6_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_3_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_62 = _tagArrayWire_6_3_T_4 | vArrayWire_6_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_7_T_1 = selArrayWire_7_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_7_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_12; // @[Cache.scala 111:28]
  wire  _tagArrayWire_7_0_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_65 = _tagArrayWire_7_0_T_4 | vArrayWire_7_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_1_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_67 = _tagArrayWire_7_1_T_4 | vArrayWire_7_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_2_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_69 = _tagArrayWire_7_2_T_4 | vArrayWire_7_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_3_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_71 = _tagArrayWire_7_3_T_4 | vArrayWire_7_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_8_T_1 = selArrayWire_8_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_8_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_14; // @[Cache.scala 111:28]
  wire  _tagArrayWire_8_0_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_74 = _tagArrayWire_8_0_T_4 | vArrayWire_8_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_1_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_76 = _tagArrayWire_8_1_T_4 | vArrayWire_8_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_2_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_78 = _tagArrayWire_8_2_T_4 | vArrayWire_8_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_3_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_80 = _tagArrayWire_8_3_T_4 | vArrayWire_8_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_9_T_1 = selArrayWire_9_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_9_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_16; // @[Cache.scala 111:28]
  wire  _tagArrayWire_9_0_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_83 = _tagArrayWire_9_0_T_4 | vArrayWire_9_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_1_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_85 = _tagArrayWire_9_1_T_4 | vArrayWire_9_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_2_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_87 = _tagArrayWire_9_2_T_4 | vArrayWire_9_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_3_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_89 = _tagArrayWire_9_3_T_4 | vArrayWire_9_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_10_T_1 = selArrayWire_10_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_10_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_18; // @[Cache.scala 111:28]
  wire  _tagArrayWire_10_0_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_92 = _tagArrayWire_10_0_T_4 | vArrayWire_10_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_1_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_94 = _tagArrayWire_10_1_T_4 | vArrayWire_10_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_2_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_96 = _tagArrayWire_10_2_T_4 | vArrayWire_10_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_3_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_98 = _tagArrayWire_10_3_T_4 | vArrayWire_10_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_11_T_1 = selArrayWire_11_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_11_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_20; // @[Cache.scala 111:28]
  wire  _tagArrayWire_11_0_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_101 = _tagArrayWire_11_0_T_4 | vArrayWire_11_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_1_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_103 = _tagArrayWire_11_1_T_4 | vArrayWire_11_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_2_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_105 = _tagArrayWire_11_2_T_4 | vArrayWire_11_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_3_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_107 = _tagArrayWire_11_3_T_4 | vArrayWire_11_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_12_T_1 = selArrayWire_12_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_12_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_22; // @[Cache.scala 111:28]
  wire  _tagArrayWire_12_0_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_110 = _tagArrayWire_12_0_T_4 | vArrayWire_12_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_1_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_112 = _tagArrayWire_12_1_T_4 | vArrayWire_12_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_2_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_114 = _tagArrayWire_12_2_T_4 | vArrayWire_12_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_3_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_116 = _tagArrayWire_12_3_T_4 | vArrayWire_12_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_13_T_1 = selArrayWire_13_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_13_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_24; // @[Cache.scala 111:28]
  wire  _tagArrayWire_13_0_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_119 = _tagArrayWire_13_0_T_4 | vArrayWire_13_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_1_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_121 = _tagArrayWire_13_1_T_4 | vArrayWire_13_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_2_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_123 = _tagArrayWire_13_2_T_4 | vArrayWire_13_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_3_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_125 = _tagArrayWire_13_3_T_4 | vArrayWire_13_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_14_T_1 = selArrayWire_14_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_14_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_26; // @[Cache.scala 111:28]
  wire  _tagArrayWire_14_0_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_128 = _tagArrayWire_14_0_T_4 | vArrayWire_14_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_1_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_130 = _tagArrayWire_14_1_T_4 | vArrayWire_14_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_2_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_132 = _tagArrayWire_14_2_T_4 | vArrayWire_14_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_3_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_134 = _tagArrayWire_14_3_T_4 | vArrayWire_14_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_15_T_1 = selArrayWire_15_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_15_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_28; // @[Cache.scala 111:28]
  wire  _tagArrayWire_15_0_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_137 = _tagArrayWire_15_0_T_4 | vArrayWire_15_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_1_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_139 = _tagArrayWire_15_1_T_4 | vArrayWire_15_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_2_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_141 = _tagArrayWire_15_2_T_4 | vArrayWire_15_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_3_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_143 = _tagArrayWire_15_3_T_4 | vArrayWire_15_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_16_T_1 = selArrayWire_16_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_16_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_30; // @[Cache.scala 111:28]
  wire  _tagArrayWire_16_0_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_146 = _tagArrayWire_16_0_T_4 | vArrayWire_16_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_1_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_148 = _tagArrayWire_16_1_T_4 | vArrayWire_16_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_2_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_150 = _tagArrayWire_16_2_T_4 | vArrayWire_16_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_3_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_152 = _tagArrayWire_16_3_T_4 | vArrayWire_16_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_17_T_1 = selArrayWire_17_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_17_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_32; // @[Cache.scala 111:28]
  wire  _tagArrayWire_17_0_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_155 = _tagArrayWire_17_0_T_4 | vArrayWire_17_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_1_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_157 = _tagArrayWire_17_1_T_4 | vArrayWire_17_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_2_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_159 = _tagArrayWire_17_2_T_4 | vArrayWire_17_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_3_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_161 = _tagArrayWire_17_3_T_4 | vArrayWire_17_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_18_T_1 = selArrayWire_18_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_18_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_34; // @[Cache.scala 111:28]
  wire  _tagArrayWire_18_0_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_164 = _tagArrayWire_18_0_T_4 | vArrayWire_18_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_1_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_166 = _tagArrayWire_18_1_T_4 | vArrayWire_18_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_2_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_168 = _tagArrayWire_18_2_T_4 | vArrayWire_18_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_3_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_170 = _tagArrayWire_18_3_T_4 | vArrayWire_18_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_19_T_1 = selArrayWire_19_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_19_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_36; // @[Cache.scala 111:28]
  wire  _tagArrayWire_19_0_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_173 = _tagArrayWire_19_0_T_4 | vArrayWire_19_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_1_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_175 = _tagArrayWire_19_1_T_4 | vArrayWire_19_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_2_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_177 = _tagArrayWire_19_2_T_4 | vArrayWire_19_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_3_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_179 = _tagArrayWire_19_3_T_4 | vArrayWire_19_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_20_T_1 = selArrayWire_20_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_20_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_38; // @[Cache.scala 111:28]
  wire  _tagArrayWire_20_0_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_182 = _tagArrayWire_20_0_T_4 | vArrayWire_20_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_1_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_184 = _tagArrayWire_20_1_T_4 | vArrayWire_20_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_2_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_186 = _tagArrayWire_20_2_T_4 | vArrayWire_20_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_3_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_188 = _tagArrayWire_20_3_T_4 | vArrayWire_20_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_21_T_1 = selArrayWire_21_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_21_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_40; // @[Cache.scala 111:28]
  wire  _tagArrayWire_21_0_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_191 = _tagArrayWire_21_0_T_4 | vArrayWire_21_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_1_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_193 = _tagArrayWire_21_1_T_4 | vArrayWire_21_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_2_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_195 = _tagArrayWire_21_2_T_4 | vArrayWire_21_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_3_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_197 = _tagArrayWire_21_3_T_4 | vArrayWire_21_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_22_T_1 = selArrayWire_22_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_22_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_42; // @[Cache.scala 111:28]
  wire  _tagArrayWire_22_0_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_200 = _tagArrayWire_22_0_T_4 | vArrayWire_22_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_1_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_202 = _tagArrayWire_22_1_T_4 | vArrayWire_22_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_2_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_204 = _tagArrayWire_22_2_T_4 | vArrayWire_22_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_3_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_206 = _tagArrayWire_22_3_T_4 | vArrayWire_22_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_23_T_1 = selArrayWire_23_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_23_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_44; // @[Cache.scala 111:28]
  wire  _tagArrayWire_23_0_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_209 = _tagArrayWire_23_0_T_4 | vArrayWire_23_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_1_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_211 = _tagArrayWire_23_1_T_4 | vArrayWire_23_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_2_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_213 = _tagArrayWire_23_2_T_4 | vArrayWire_23_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_3_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_215 = _tagArrayWire_23_3_T_4 | vArrayWire_23_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_24_T_1 = selArrayWire_24_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_24_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_46; // @[Cache.scala 111:28]
  wire  _tagArrayWire_24_0_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_218 = _tagArrayWire_24_0_T_4 | vArrayWire_24_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_1_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_220 = _tagArrayWire_24_1_T_4 | vArrayWire_24_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_2_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_222 = _tagArrayWire_24_2_T_4 | vArrayWire_24_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_3_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_224 = _tagArrayWire_24_3_T_4 | vArrayWire_24_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_25_T_1 = selArrayWire_25_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_25_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_48; // @[Cache.scala 111:28]
  wire  _tagArrayWire_25_0_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_227 = _tagArrayWire_25_0_T_4 | vArrayWire_25_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_1_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_229 = _tagArrayWire_25_1_T_4 | vArrayWire_25_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_2_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_231 = _tagArrayWire_25_2_T_4 | vArrayWire_25_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_3_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_233 = _tagArrayWire_25_3_T_4 | vArrayWire_25_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_26_T_1 = selArrayWire_26_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_26_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_50; // @[Cache.scala 111:28]
  wire  _tagArrayWire_26_0_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_236 = _tagArrayWire_26_0_T_4 | vArrayWire_26_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_1_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_238 = _tagArrayWire_26_1_T_4 | vArrayWire_26_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_2_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_240 = _tagArrayWire_26_2_T_4 | vArrayWire_26_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_3_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_242 = _tagArrayWire_26_3_T_4 | vArrayWire_26_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_27_T_1 = selArrayWire_27_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_27_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_52; // @[Cache.scala 111:28]
  wire  _tagArrayWire_27_0_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_245 = _tagArrayWire_27_0_T_4 | vArrayWire_27_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_1_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_247 = _tagArrayWire_27_1_T_4 | vArrayWire_27_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_2_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_249 = _tagArrayWire_27_2_T_4 | vArrayWire_27_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_3_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_251 = _tagArrayWire_27_3_T_4 | vArrayWire_27_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_28_T_1 = selArrayWire_28_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_28_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_54; // @[Cache.scala 111:28]
  wire  _tagArrayWire_28_0_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_254 = _tagArrayWire_28_0_T_4 | vArrayWire_28_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_1_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_256 = _tagArrayWire_28_1_T_4 | vArrayWire_28_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_2_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_258 = _tagArrayWire_28_2_T_4 | vArrayWire_28_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_3_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_260 = _tagArrayWire_28_3_T_4 | vArrayWire_28_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_29_T_1 = selArrayWire_29_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_29_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_56; // @[Cache.scala 111:28]
  wire  _tagArrayWire_29_0_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_263 = _tagArrayWire_29_0_T_4 | vArrayWire_29_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_1_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_265 = _tagArrayWire_29_1_T_4 | vArrayWire_29_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_2_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_267 = _tagArrayWire_29_2_T_4 | vArrayWire_29_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_3_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_269 = _tagArrayWire_29_3_T_4 | vArrayWire_29_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_30_T_1 = selArrayWire_30_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_30_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_58; // @[Cache.scala 111:28]
  wire  _tagArrayWire_30_0_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_272 = _tagArrayWire_30_0_T_4 | vArrayWire_30_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_1_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_274 = _tagArrayWire_30_1_T_4 | vArrayWire_30_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_2_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_276 = _tagArrayWire_30_2_T_4 | vArrayWire_30_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_3_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_278 = _tagArrayWire_30_3_T_4 | vArrayWire_30_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_31_T_1 = selArrayWire_31_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_31_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_60; // @[Cache.scala 111:28]
  wire  _tagArrayWire_31_0_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_281 = _tagArrayWire_31_0_T_4 | vArrayWire_31_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_1_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_283 = _tagArrayWire_31_1_T_4 | vArrayWire_31_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_2_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_285 = _tagArrayWire_31_2_T_4 | vArrayWire_31_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_3_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_287 = _tagArrayWire_31_3_T_4 | vArrayWire_31_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_32_T_1 = selArrayWire_32_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_32_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_62; // @[Cache.scala 111:28]
  wire  _tagArrayWire_32_0_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_290 = _tagArrayWire_32_0_T_4 | vArrayWire_32_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_1_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_292 = _tagArrayWire_32_1_T_4 | vArrayWire_32_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_2_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_294 = _tagArrayWire_32_2_T_4 | vArrayWire_32_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_3_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_296 = _tagArrayWire_32_3_T_4 | vArrayWire_32_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_33_T_1 = selArrayWire_33_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_33_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_64; // @[Cache.scala 111:28]
  wire  _tagArrayWire_33_0_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_299 = _tagArrayWire_33_0_T_4 | vArrayWire_33_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_1_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_301 = _tagArrayWire_33_1_T_4 | vArrayWire_33_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_2_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_303 = _tagArrayWire_33_2_T_4 | vArrayWire_33_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_3_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_305 = _tagArrayWire_33_3_T_4 | vArrayWire_33_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_34_T_1 = selArrayWire_34_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_34_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_66; // @[Cache.scala 111:28]
  wire  _tagArrayWire_34_0_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_308 = _tagArrayWire_34_0_T_4 | vArrayWire_34_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_1_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_310 = _tagArrayWire_34_1_T_4 | vArrayWire_34_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_2_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_312 = _tagArrayWire_34_2_T_4 | vArrayWire_34_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_3_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_314 = _tagArrayWire_34_3_T_4 | vArrayWire_34_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_35_T_1 = selArrayWire_35_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_35_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_68; // @[Cache.scala 111:28]
  wire  _tagArrayWire_35_0_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_317 = _tagArrayWire_35_0_T_4 | vArrayWire_35_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_1_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_319 = _tagArrayWire_35_1_T_4 | vArrayWire_35_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_2_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_321 = _tagArrayWire_35_2_T_4 | vArrayWire_35_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_3_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_323 = _tagArrayWire_35_3_T_4 | vArrayWire_35_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_36_T_1 = selArrayWire_36_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_36_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_70; // @[Cache.scala 111:28]
  wire  _tagArrayWire_36_0_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_326 = _tagArrayWire_36_0_T_4 | vArrayWire_36_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_1_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_328 = _tagArrayWire_36_1_T_4 | vArrayWire_36_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_2_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_330 = _tagArrayWire_36_2_T_4 | vArrayWire_36_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_3_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_332 = _tagArrayWire_36_3_T_4 | vArrayWire_36_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_37_T_1 = selArrayWire_37_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_37_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_72; // @[Cache.scala 111:28]
  wire  _tagArrayWire_37_0_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_335 = _tagArrayWire_37_0_T_4 | vArrayWire_37_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_1_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_337 = _tagArrayWire_37_1_T_4 | vArrayWire_37_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_2_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_339 = _tagArrayWire_37_2_T_4 | vArrayWire_37_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_3_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_341 = _tagArrayWire_37_3_T_4 | vArrayWire_37_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_38_T_1 = selArrayWire_38_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_38_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_74; // @[Cache.scala 111:28]
  wire  _tagArrayWire_38_0_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_344 = _tagArrayWire_38_0_T_4 | vArrayWire_38_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_1_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_346 = _tagArrayWire_38_1_T_4 | vArrayWire_38_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_2_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_348 = _tagArrayWire_38_2_T_4 | vArrayWire_38_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_3_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_350 = _tagArrayWire_38_3_T_4 | vArrayWire_38_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_39_T_1 = selArrayWire_39_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_39_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_76; // @[Cache.scala 111:28]
  wire  _tagArrayWire_39_0_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_353 = _tagArrayWire_39_0_T_4 | vArrayWire_39_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_1_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_355 = _tagArrayWire_39_1_T_4 | vArrayWire_39_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_2_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_357 = _tagArrayWire_39_2_T_4 | vArrayWire_39_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_3_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_359 = _tagArrayWire_39_3_T_4 | vArrayWire_39_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_40_T_1 = selArrayWire_40_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_40_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_78; // @[Cache.scala 111:28]
  wire  _tagArrayWire_40_0_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_362 = _tagArrayWire_40_0_T_4 | vArrayWire_40_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_1_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_364 = _tagArrayWire_40_1_T_4 | vArrayWire_40_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_2_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_366 = _tagArrayWire_40_2_T_4 | vArrayWire_40_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_3_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_368 = _tagArrayWire_40_3_T_4 | vArrayWire_40_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_41_T_1 = selArrayWire_41_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_41_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_80; // @[Cache.scala 111:28]
  wire  _tagArrayWire_41_0_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_371 = _tagArrayWire_41_0_T_4 | vArrayWire_41_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_1_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_373 = _tagArrayWire_41_1_T_4 | vArrayWire_41_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_2_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_375 = _tagArrayWire_41_2_T_4 | vArrayWire_41_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_3_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_377 = _tagArrayWire_41_3_T_4 | vArrayWire_41_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_42_T_1 = selArrayWire_42_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_42_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_82; // @[Cache.scala 111:28]
  wire  _tagArrayWire_42_0_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_380 = _tagArrayWire_42_0_T_4 | vArrayWire_42_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_1_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_382 = _tagArrayWire_42_1_T_4 | vArrayWire_42_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_2_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_384 = _tagArrayWire_42_2_T_4 | vArrayWire_42_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_3_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_386 = _tagArrayWire_42_3_T_4 | vArrayWire_42_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_43_T_1 = selArrayWire_43_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_43_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_84; // @[Cache.scala 111:28]
  wire  _tagArrayWire_43_0_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_389 = _tagArrayWire_43_0_T_4 | vArrayWire_43_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_1_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_391 = _tagArrayWire_43_1_T_4 | vArrayWire_43_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_2_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_393 = _tagArrayWire_43_2_T_4 | vArrayWire_43_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_3_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_395 = _tagArrayWire_43_3_T_4 | vArrayWire_43_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_44_T_1 = selArrayWire_44_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_44_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_86; // @[Cache.scala 111:28]
  wire  _tagArrayWire_44_0_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_398 = _tagArrayWire_44_0_T_4 | vArrayWire_44_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_1_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_400 = _tagArrayWire_44_1_T_4 | vArrayWire_44_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_2_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_402 = _tagArrayWire_44_2_T_4 | vArrayWire_44_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_3_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_404 = _tagArrayWire_44_3_T_4 | vArrayWire_44_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_45_T_1 = selArrayWire_45_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_45_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_88; // @[Cache.scala 111:28]
  wire  _tagArrayWire_45_0_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_407 = _tagArrayWire_45_0_T_4 | vArrayWire_45_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_1_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_409 = _tagArrayWire_45_1_T_4 | vArrayWire_45_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_2_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_411 = _tagArrayWire_45_2_T_4 | vArrayWire_45_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_3_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_413 = _tagArrayWire_45_3_T_4 | vArrayWire_45_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_46_T_1 = selArrayWire_46_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_46_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_90; // @[Cache.scala 111:28]
  wire  _tagArrayWire_46_0_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_416 = _tagArrayWire_46_0_T_4 | vArrayWire_46_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_1_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_418 = _tagArrayWire_46_1_T_4 | vArrayWire_46_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_2_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_420 = _tagArrayWire_46_2_T_4 | vArrayWire_46_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_3_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_422 = _tagArrayWire_46_3_T_4 | vArrayWire_46_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_47_T_1 = selArrayWire_47_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_47_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_92; // @[Cache.scala 111:28]
  wire  _tagArrayWire_47_0_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_425 = _tagArrayWire_47_0_T_4 | vArrayWire_47_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_1_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_427 = _tagArrayWire_47_1_T_4 | vArrayWire_47_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_2_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_429 = _tagArrayWire_47_2_T_4 | vArrayWire_47_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_3_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_431 = _tagArrayWire_47_3_T_4 | vArrayWire_47_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_48_T_1 = selArrayWire_48_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_48_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_94; // @[Cache.scala 111:28]
  wire  _tagArrayWire_48_0_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_434 = _tagArrayWire_48_0_T_4 | vArrayWire_48_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_1_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_436 = _tagArrayWire_48_1_T_4 | vArrayWire_48_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_2_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_438 = _tagArrayWire_48_2_T_4 | vArrayWire_48_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_3_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_440 = _tagArrayWire_48_3_T_4 | vArrayWire_48_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_49_T_1 = selArrayWire_49_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_49_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_96; // @[Cache.scala 111:28]
  wire  _tagArrayWire_49_0_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_443 = _tagArrayWire_49_0_T_4 | vArrayWire_49_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_1_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_445 = _tagArrayWire_49_1_T_4 | vArrayWire_49_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_2_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_447 = _tagArrayWire_49_2_T_4 | vArrayWire_49_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_3_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_449 = _tagArrayWire_49_3_T_4 | vArrayWire_49_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_50_T_1 = selArrayWire_50_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_50_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_98; // @[Cache.scala 111:28]
  wire  _tagArrayWire_50_0_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_452 = _tagArrayWire_50_0_T_4 | vArrayWire_50_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_1_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_454 = _tagArrayWire_50_1_T_4 | vArrayWire_50_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_2_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_456 = _tagArrayWire_50_2_T_4 | vArrayWire_50_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_3_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_458 = _tagArrayWire_50_3_T_4 | vArrayWire_50_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_51_T_1 = selArrayWire_51_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_51_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_100; // @[Cache.scala 111:28]
  wire  _tagArrayWire_51_0_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_461 = _tagArrayWire_51_0_T_4 | vArrayWire_51_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_1_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_463 = _tagArrayWire_51_1_T_4 | vArrayWire_51_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_2_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_465 = _tagArrayWire_51_2_T_4 | vArrayWire_51_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_3_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_467 = _tagArrayWire_51_3_T_4 | vArrayWire_51_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_52_T_1 = selArrayWire_52_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_52_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_102; // @[Cache.scala 111:28]
  wire  _tagArrayWire_52_0_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_470 = _tagArrayWire_52_0_T_4 | vArrayWire_52_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_1_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_472 = _tagArrayWire_52_1_T_4 | vArrayWire_52_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_2_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_474 = _tagArrayWire_52_2_T_4 | vArrayWire_52_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_3_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_476 = _tagArrayWire_52_3_T_4 | vArrayWire_52_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_53_T_1 = selArrayWire_53_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_53_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_104; // @[Cache.scala 111:28]
  wire  _tagArrayWire_53_0_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_479 = _tagArrayWire_53_0_T_4 | vArrayWire_53_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_1_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_481 = _tagArrayWire_53_1_T_4 | vArrayWire_53_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_2_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_483 = _tagArrayWire_53_2_T_4 | vArrayWire_53_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_3_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_485 = _tagArrayWire_53_3_T_4 | vArrayWire_53_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_54_T_1 = selArrayWire_54_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_54_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_106; // @[Cache.scala 111:28]
  wire  _tagArrayWire_54_0_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_488 = _tagArrayWire_54_0_T_4 | vArrayWire_54_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_1_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_490 = _tagArrayWire_54_1_T_4 | vArrayWire_54_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_2_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_492 = _tagArrayWire_54_2_T_4 | vArrayWire_54_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_3_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_494 = _tagArrayWire_54_3_T_4 | vArrayWire_54_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_55_T_1 = selArrayWire_55_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_55_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_108; // @[Cache.scala 111:28]
  wire  _tagArrayWire_55_0_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_497 = _tagArrayWire_55_0_T_4 | vArrayWire_55_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_1_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_499 = _tagArrayWire_55_1_T_4 | vArrayWire_55_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_2_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_501 = _tagArrayWire_55_2_T_4 | vArrayWire_55_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_3_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_503 = _tagArrayWire_55_3_T_4 | vArrayWire_55_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_56_T_1 = selArrayWire_56_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_56_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_110; // @[Cache.scala 111:28]
  wire  _tagArrayWire_56_0_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_506 = _tagArrayWire_56_0_T_4 | vArrayWire_56_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_1_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_508 = _tagArrayWire_56_1_T_4 | vArrayWire_56_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_2_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_510 = _tagArrayWire_56_2_T_4 | vArrayWire_56_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_3_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_512 = _tagArrayWire_56_3_T_4 | vArrayWire_56_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_57_T_1 = selArrayWire_57_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_57_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_112; // @[Cache.scala 111:28]
  wire  _tagArrayWire_57_0_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_515 = _tagArrayWire_57_0_T_4 | vArrayWire_57_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_1_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_517 = _tagArrayWire_57_1_T_4 | vArrayWire_57_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_2_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_519 = _tagArrayWire_57_2_T_4 | vArrayWire_57_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_3_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_521 = _tagArrayWire_57_3_T_4 | vArrayWire_57_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_58_T_1 = selArrayWire_58_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_58_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_114; // @[Cache.scala 111:28]
  wire  _tagArrayWire_58_0_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_524 = _tagArrayWire_58_0_T_4 | vArrayWire_58_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_1_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_526 = _tagArrayWire_58_1_T_4 | vArrayWire_58_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_2_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_528 = _tagArrayWire_58_2_T_4 | vArrayWire_58_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_3_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_530 = _tagArrayWire_58_3_T_4 | vArrayWire_58_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_59_T_1 = selArrayWire_59_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_59_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_116; // @[Cache.scala 111:28]
  wire  _tagArrayWire_59_0_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_533 = _tagArrayWire_59_0_T_4 | vArrayWire_59_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_1_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_535 = _tagArrayWire_59_1_T_4 | vArrayWire_59_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_2_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_537 = _tagArrayWire_59_2_T_4 | vArrayWire_59_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_3_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_539 = _tagArrayWire_59_3_T_4 | vArrayWire_59_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_60_T_1 = selArrayWire_60_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_60_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_118; // @[Cache.scala 111:28]
  wire  _tagArrayWire_60_0_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_542 = _tagArrayWire_60_0_T_4 | vArrayWire_60_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_1_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_544 = _tagArrayWire_60_1_T_4 | vArrayWire_60_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_2_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_546 = _tagArrayWire_60_2_T_4 | vArrayWire_60_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_3_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_548 = _tagArrayWire_60_3_T_4 | vArrayWire_60_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_61_T_1 = selArrayWire_61_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_61_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_120; // @[Cache.scala 111:28]
  wire  _tagArrayWire_61_0_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_551 = _tagArrayWire_61_0_T_4 | vArrayWire_61_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_1_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_553 = _tagArrayWire_61_1_T_4 | vArrayWire_61_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_2_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_555 = _tagArrayWire_61_2_T_4 | vArrayWire_61_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_3_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_557 = _tagArrayWire_61_3_T_4 | vArrayWire_61_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_62_T_1 = selArrayWire_62_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_62_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_122; // @[Cache.scala 111:28]
  wire  _tagArrayWire_62_0_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_560 = _tagArrayWire_62_0_T_4 | vArrayWire_62_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_1_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_562 = _tagArrayWire_62_1_T_4 | vArrayWire_62_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_2_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_564 = _tagArrayWire_62_2_T_4 | vArrayWire_62_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_3_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_566 = _tagArrayWire_62_3_T_4 | vArrayWire_62_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_63_T_1 = selArrayWire_63_r + 2'h1; // @[Cache.scala 109:23]
  wire  _selArrayWire_63_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_124; // @[Cache.scala 111:28]
  wire  _tagArrayWire_63_0_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h0 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_569 = _tagArrayWire_63_0_T_4 | vArrayWire_63_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_1_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h1 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_571 = _tagArrayWire_63_1_T_4 | vArrayWire_63_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_2_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h2 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_573 = _tagArrayWire_63_2_T_4 | vArrayWire_63_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_3_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h3 & cacheState; // @[Cache.scala 114:112]
  wire  _GEN_575 = _tagArrayWire_63_3_T_4 | vArrayWire_63_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _io_SRAMIO_0_cen_T_2 = cacheState & io_cacheOut_r_valid_i & 2'h0 == sramSel; // @[Cache.scala 147:52]
  wire [127:0] _io_SRAMIO_0_wdata_T = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _io_SRAMIO_0_wdata_T_1 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 30:58]
  wire  _io_SRAMIO_1_cen_T_2 = cacheState & io_cacheOut_r_valid_i & 2'h1 == sramSel; // @[Cache.scala 147:52]
  wire  _io_SRAMIO_2_cen_T_2 = cacheState & io_cacheOut_r_valid_i & 2'h2 == sramSel; // @[Cache.scala 147:52]
  wire  _io_SRAMIO_3_cen_T_2 = cacheState & io_cacheOut_r_valid_i & 2'h3 == sramSel; // @[Cache.scala 147:52]
  assign io_cacheOut_ar_valid_o = cacheState; // @[Cache.scala 46:27]
  assign io_cacheOut_ar_addr_o = {io_cacheOut_ar_addr_o_hi,4'h0}; // @[Cat.scala 30:58]
  assign io_cacheOut_ar_len_o = {{7'd0}, cacheState}; // @[Cache.scala 46:27]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 139:24]
  assign io_cacheIn_ready = isIdle & hit; // @[Cache.scala 155:30]
  assign io_cacheIn_data_read = offset[3] ? waysel[127:64] : waysel[63:0]; // @[Cache.scala 92:30]
  assign io_SRAMIO_0_cen = ~(cacheState & io_cacheOut_r_valid_i & 2'h0 == sramSel); // @[Cache.scala 147:16]
  assign io_SRAMIO_0_wen = ~_io_SRAMIO_0_cen_T_2; // @[Cache.scala 149:16]
  assign io_SRAMIO_0_wdata = io_cacheOut_r_last_i ? _io_SRAMIO_0_wdata_T : _io_SRAMIO_0_wdata_T_1; // @[Cache.scala 150:21]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  assign io_SRAMIO_0_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:21]
  assign io_SRAMIO_1_cen = ~(cacheState & io_cacheOut_r_valid_i & 2'h1 == sramSel); // @[Cache.scala 147:16]
  assign io_SRAMIO_1_wen = ~_io_SRAMIO_1_cen_T_2; // @[Cache.scala 149:16]
  assign io_SRAMIO_1_wdata = io_cacheOut_r_last_i ? _io_SRAMIO_0_wdata_T : _io_SRAMIO_0_wdata_T_1; // @[Cache.scala 150:21]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  assign io_SRAMIO_1_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:21]
  assign io_SRAMIO_2_cen = ~(cacheState & io_cacheOut_r_valid_i & 2'h2 == sramSel); // @[Cache.scala 147:16]
  assign io_SRAMIO_2_wen = ~_io_SRAMIO_2_cen_T_2; // @[Cache.scala 149:16]
  assign io_SRAMIO_2_wdata = io_cacheOut_r_last_i ? _io_SRAMIO_0_wdata_T : _io_SRAMIO_0_wdata_T_1; // @[Cache.scala 150:21]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  assign io_SRAMIO_2_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:21]
  assign io_SRAMIO_3_cen = ~(cacheState & io_cacheOut_r_valid_i & 2'h3 == sramSel); // @[Cache.scala 147:16]
  assign io_SRAMIO_3_wen = ~_io_SRAMIO_3_cen_T_2; // @[Cache.scala 149:16]
  assign io_SRAMIO_3_wdata = io_cacheOut_r_last_i ? _io_SRAMIO_0_wdata_T : _io_SRAMIO_0_wdata_T_1; // @[Cache.scala 150:21]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 28:30]
  assign io_SRAMIO_3_wmask = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000; // @[Cache.scala 151:21]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 32:27]
      cacheState <= 1'h0; // @[Cache.scala 32:27]
    end else if (cacheState) begin // @[Mux.scala 80:57]
      if (io_cacheOut_r_last_i) begin // @[Cache.scala 36:20]
        cacheState <= 1'h0;
      end else begin
        cacheState <= 1'h1;
      end
    end else begin
      cacheState <= IdleMux;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_63_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_0_r <= _GEN_569;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_62_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_0_r <= _GEN_560;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_61_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_0_r <= _GEN_551;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_60_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_0_r <= _GEN_542;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_59_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_0_r <= _GEN_533;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_58_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_0_r <= _GEN_524;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_57_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_0_r <= _GEN_515;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_56_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_0_r <= _GEN_506;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_55_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_0_r <= _GEN_497;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_54_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_0_r <= _GEN_488;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_53_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_0_r <= _GEN_479;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_52_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_0_r <= _GEN_470;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_51_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_0_r <= _GEN_461;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_50_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_0_r <= _GEN_452;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_49_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_0_r <= _GEN_443;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_48_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_0_r <= _GEN_434;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_47_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_0_r <= _GEN_425;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_46_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_0_r <= _GEN_416;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_45_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_0_r <= _GEN_407;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_44_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_0_r <= _GEN_398;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_43_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_0_r <= _GEN_389;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_42_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_0_r <= _GEN_380;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_41_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_0_r <= _GEN_371;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_40_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_0_r <= _GEN_362;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_39_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_0_r <= _GEN_353;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_38_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_0_r <= _GEN_344;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_37_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_0_r <= _GEN_335;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_36_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_0_r <= _GEN_326;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_35_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_0_r <= _GEN_317;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_34_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_0_r <= _GEN_308;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_33_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_0_r <= _GEN_299;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_32_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_0_r <= _GEN_290;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_31_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_0_r <= _GEN_281;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_30_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_0_r <= _GEN_272;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_29_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_0_r <= _GEN_263;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_28_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_0_r <= _GEN_254;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_27_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_0_r <= _GEN_245;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_26_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_0_r <= _GEN_236;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_25_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_0_r <= _GEN_227;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_24_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_0_r <= _GEN_218;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_23_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_0_r <= _GEN_209;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_22_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_0_r <= _GEN_200;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_21_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_0_r <= _GEN_191;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_20_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_0_r <= _GEN_182;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_19_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_0_r <= _GEN_173;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_18_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_0_r <= _GEN_164;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_17_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_0_r <= _GEN_155;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_16_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_0_r <= _GEN_146;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_15_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_0_r <= _GEN_137;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_14_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_0_r <= _GEN_128;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_13_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_0_r <= _GEN_119;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_12_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_0_r <= _GEN_110;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_11_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_0_r <= _GEN_101;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_10_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_0_r <= _GEN_92;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_9_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_0_r <= _GEN_83;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_8_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_0_r <= _GEN_74;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_7_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_0_r <= _GEN_65;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_6_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_0_r <= _GEN_56;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_5_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_0_r <= _GEN_47;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_4_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_0_r <= _GEN_38;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_3_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_0_r <= _GEN_29;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_2_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_0_r <= _GEN_20;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_1_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_0_r <= _GEN_11;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_0_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_0_r <= _GEN_2;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_63_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_1_r <= _GEN_571;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_62_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_1_r <= _GEN_562;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_61_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_1_r <= _GEN_553;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_60_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_1_r <= _GEN_544;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_59_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_1_r <= _GEN_535;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_58_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_1_r <= _GEN_526;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_57_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_1_r <= _GEN_517;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_56_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_1_r <= _GEN_508;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_55_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_1_r <= _GEN_499;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_54_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_1_r <= _GEN_490;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_53_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_1_r <= _GEN_481;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_52_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_1_r <= _GEN_472;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_51_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_1_r <= _GEN_463;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_50_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_1_r <= _GEN_454;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_49_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_1_r <= _GEN_445;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_48_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_1_r <= _GEN_436;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_47_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_1_r <= _GEN_427;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_46_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_1_r <= _GEN_418;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_45_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_1_r <= _GEN_409;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_44_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_1_r <= _GEN_400;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_43_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_1_r <= _GEN_391;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_42_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_1_r <= _GEN_382;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_41_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_1_r <= _GEN_373;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_40_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_1_r <= _GEN_364;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_39_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_1_r <= _GEN_355;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_38_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_1_r <= _GEN_346;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_37_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_1_r <= _GEN_337;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_36_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_1_r <= _GEN_328;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_35_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_1_r <= _GEN_319;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_34_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_1_r <= _GEN_310;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_33_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_1_r <= _GEN_301;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_32_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_1_r <= _GEN_292;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_31_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_1_r <= _GEN_283;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_30_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_1_r <= _GEN_274;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_29_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_1_r <= _GEN_265;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_28_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_1_r <= _GEN_256;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_27_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_1_r <= _GEN_247;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_26_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_1_r <= _GEN_238;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_25_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_1_r <= _GEN_229;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_24_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_1_r <= _GEN_220;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_23_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_1_r <= _GEN_211;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_22_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_1_r <= _GEN_202;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_21_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_1_r <= _GEN_193;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_20_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_1_r <= _GEN_184;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_19_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_1_r <= _GEN_175;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_18_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_1_r <= _GEN_166;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_17_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_1_r <= _GEN_157;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_16_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_1_r <= _GEN_148;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_15_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_1_r <= _GEN_139;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_14_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_1_r <= _GEN_130;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_13_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_1_r <= _GEN_121;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_12_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_1_r <= _GEN_112;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_11_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_1_r <= _GEN_103;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_10_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_1_r <= _GEN_94;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_9_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_1_r <= _GEN_85;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_8_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_1_r <= _GEN_76;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_7_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_1_r <= _GEN_67;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_6_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_1_r <= _GEN_58;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_5_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_1_r <= _GEN_49;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_4_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_1_r <= _GEN_40;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_3_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_1_r <= _GEN_31;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_2_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_1_r <= _GEN_22;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_1_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_1_r <= _GEN_13;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_0_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_1_r <= _GEN_4;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_63_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_2_r <= _GEN_573;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_62_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_2_r <= _GEN_564;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_61_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_2_r <= _GEN_555;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_60_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_2_r <= _GEN_546;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_59_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_2_r <= _GEN_537;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_58_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_2_r <= _GEN_528;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_57_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_2_r <= _GEN_519;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_56_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_2_r <= _GEN_510;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_55_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_2_r <= _GEN_501;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_54_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_2_r <= _GEN_492;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_53_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_2_r <= _GEN_483;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_52_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_2_r <= _GEN_474;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_51_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_2_r <= _GEN_465;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_50_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_2_r <= _GEN_456;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_49_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_2_r <= _GEN_447;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_48_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_2_r <= _GEN_438;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_47_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_2_r <= _GEN_429;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_46_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_2_r <= _GEN_420;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_45_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_2_r <= _GEN_411;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_44_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_2_r <= _GEN_402;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_43_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_2_r <= _GEN_393;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_42_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_2_r <= _GEN_384;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_41_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_2_r <= _GEN_375;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_40_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_2_r <= _GEN_366;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_39_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_2_r <= _GEN_357;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_38_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_2_r <= _GEN_348;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_37_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_2_r <= _GEN_339;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_36_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_2_r <= _GEN_330;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_35_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_2_r <= _GEN_321;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_34_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_2_r <= _GEN_312;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_33_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_2_r <= _GEN_303;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_32_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_2_r <= _GEN_294;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_31_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_2_r <= _GEN_285;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_30_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_2_r <= _GEN_276;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_29_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_2_r <= _GEN_267;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_28_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_2_r <= _GEN_258;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_27_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_2_r <= _GEN_249;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_26_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_2_r <= _GEN_240;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_25_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_2_r <= _GEN_231;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_24_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_2_r <= _GEN_222;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_23_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_2_r <= _GEN_213;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_22_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_2_r <= _GEN_204;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_21_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_2_r <= _GEN_195;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_20_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_2_r <= _GEN_186;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_19_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_2_r <= _GEN_177;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_18_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_2_r <= _GEN_168;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_17_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_2_r <= _GEN_159;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_16_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_2_r <= _GEN_150;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_15_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_2_r <= _GEN_141;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_14_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_2_r <= _GEN_132;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_13_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_2_r <= _GEN_123;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_12_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_2_r <= _GEN_114;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_11_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_2_r <= _GEN_105;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_10_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_2_r <= _GEN_96;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_9_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_2_r <= _GEN_87;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_8_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_2_r <= _GEN_78;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_7_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_2_r <= _GEN_69;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_6_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_2_r <= _GEN_60;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_5_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_2_r <= _GEN_51;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_4_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_2_r <= _GEN_42;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_3_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_2_r <= _GEN_33;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_2_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_2_r <= _GEN_24;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_1_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_2_r <= _GEN_15;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_0_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_2_r <= _GEN_6;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_63_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_3_r <= _GEN_575;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_62_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_3_r <= _GEN_566;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_61_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_3_r <= _GEN_557;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_60_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_3_r <= _GEN_548;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_59_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_3_r <= _GEN_539;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_58_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_3_r <= _GEN_530;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_57_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_3_r <= _GEN_521;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_56_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_3_r <= _GEN_512;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_55_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_3_r <= _GEN_503;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_54_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_3_r <= _GEN_494;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_53_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_3_r <= _GEN_485;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_52_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_3_r <= _GEN_476;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_51_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_3_r <= _GEN_467;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_50_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_3_r <= _GEN_458;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_49_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_3_r <= _GEN_449;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_48_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_3_r <= _GEN_440;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_47_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_3_r <= _GEN_431;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_46_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_3_r <= _GEN_422;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_45_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_3_r <= _GEN_413;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_44_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_3_r <= _GEN_404;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_43_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_3_r <= _GEN_395;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_42_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_3_r <= _GEN_386;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_41_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_3_r <= _GEN_377;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_40_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_3_r <= _GEN_368;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_39_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_3_r <= _GEN_359;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_38_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_3_r <= _GEN_350;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_37_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_3_r <= _GEN_341;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_36_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_3_r <= _GEN_332;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_35_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_3_r <= _GEN_323;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_34_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_3_r <= _GEN_314;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_33_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_3_r <= _GEN_305;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_32_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_3_r <= _GEN_296;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_31_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_3_r <= _GEN_287;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_30_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_3_r <= _GEN_278;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_29_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_3_r <= _GEN_269;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_28_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_3_r <= _GEN_260;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_27_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_3_r <= _GEN_251;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_26_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_3_r <= _GEN_242;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_25_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_3_r <= _GEN_233;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_24_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_3_r <= _GEN_224;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_23_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_3_r <= _GEN_215;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_22_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_3_r <= _GEN_206;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_21_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_3_r <= _GEN_197;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_20_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_3_r <= _GEN_188;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_19_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_3_r <= _GEN_179;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_18_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_3_r <= _GEN_170;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_17_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_3_r <= _GEN_161;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_16_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_3_r <= _GEN_152;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_15_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_3_r <= _GEN_143;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_14_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_3_r <= _GEN_134;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_13_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_3_r <= _GEN_125;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_12_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_3_r <= _GEN_116;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_11_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_3_r <= _GEN_107;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_10_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_3_r <= _GEN_98;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_9_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_3_r <= _GEN_89;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_8_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_3_r <= _GEN_80;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_7_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_3_r <= _GEN_71;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_6_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_3_r <= _GEN_62;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_5_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_3_r <= _GEN_53;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_4_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_3_r <= _GEN_44;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_3_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_3_r <= _GEN_35;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_2_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_3_r <= _GEN_26;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_1_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_3_r <= _GEN_17;
    end
    if (_T_1) begin // @[Reg.scala 27:20]
      vArrayWire_0_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_3_r <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_1_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_1_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_1_r <= _selArrayWire_1_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_0_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_0_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_0_r <= _selArrayWire_0_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_2_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_2_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_2_r <= _selArrayWire_2_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_3_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_3_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_3_r <= _selArrayWire_3_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_4_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_4_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_4_r <= _selArrayWire_4_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_5_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_5_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_5_r <= _selArrayWire_5_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_6_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_6_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_6_r <= _selArrayWire_6_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_7_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_7_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_7_r <= _selArrayWire_7_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_8_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_8_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_8_r <= _selArrayWire_8_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_9_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_9_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_9_r <= _selArrayWire_9_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_10_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_10_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_10_r <= _selArrayWire_10_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_11_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_11_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_11_r <= _selArrayWire_11_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_12_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_12_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_12_r <= _selArrayWire_12_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_13_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_13_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_13_r <= _selArrayWire_13_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_14_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_14_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_14_r <= _selArrayWire_14_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_15_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_15_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_15_r <= _selArrayWire_15_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_16_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_16_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_16_r <= _selArrayWire_16_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_17_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_17_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_17_r <= _selArrayWire_17_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_18_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_18_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_18_r <= _selArrayWire_18_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_19_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_19_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_19_r <= _selArrayWire_19_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_20_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_20_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_20_r <= _selArrayWire_20_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_21_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_21_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_21_r <= _selArrayWire_21_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_22_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_22_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_22_r <= _selArrayWire_22_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_23_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_23_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_23_r <= _selArrayWire_23_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_24_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_24_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_24_r <= _selArrayWire_24_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_25_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_25_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_25_r <= _selArrayWire_25_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_26_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_26_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_26_r <= _selArrayWire_26_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_27_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_27_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_27_r <= _selArrayWire_27_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_28_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_28_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_28_r <= _selArrayWire_28_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_29_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_29_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_29_r <= _selArrayWire_29_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_30_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_30_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_30_r <= _selArrayWire_30_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_31_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_31_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_31_r <= _selArrayWire_31_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_32_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_32_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_32_r <= _selArrayWire_32_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_33_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_33_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_33_r <= _selArrayWire_33_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_34_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_34_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_34_r <= _selArrayWire_34_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_35_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_35_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_35_r <= _selArrayWire_35_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_36_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_36_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_36_r <= _selArrayWire_36_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_37_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_37_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_37_r <= _selArrayWire_37_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_38_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_38_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_38_r <= _selArrayWire_38_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_39_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_39_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_39_r <= _selArrayWire_39_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_40_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_40_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_40_r <= _selArrayWire_40_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_41_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_41_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_41_r <= _selArrayWire_41_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_42_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_42_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_42_r <= _selArrayWire_42_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_43_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_43_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_43_r <= _selArrayWire_43_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_44_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_44_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_44_r <= _selArrayWire_44_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_45_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_45_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_45_r <= _selArrayWire_45_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_46_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_46_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_46_r <= _selArrayWire_46_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_47_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_47_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_47_r <= _selArrayWire_47_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_48_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_48_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_48_r <= _selArrayWire_48_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_49_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_49_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_49_r <= _selArrayWire_49_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_50_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_50_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_50_r <= _selArrayWire_50_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_51_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_51_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_51_r <= _selArrayWire_51_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_52_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_52_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_52_r <= _selArrayWire_52_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_53_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_53_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_53_r <= _selArrayWire_53_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_54_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_54_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_54_r <= _selArrayWire_54_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_55_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_55_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_55_r <= _selArrayWire_55_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_56_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_56_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_56_r <= _selArrayWire_56_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_57_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_57_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_57_r <= _selArrayWire_57_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_58_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_58_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_58_r <= _selArrayWire_58_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_59_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_59_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_59_r <= _selArrayWire_59_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_60_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_60_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_60_r <= _selArrayWire_60_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_61_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_61_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_61_r <= _selArrayWire_61_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_62_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_62_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_62_r <= _selArrayWire_62_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_63_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_63_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_63_r <= _selArrayWire_63_T_1; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cacheState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  vArrayWire_63_0_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vArrayWire_62_0_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  vArrayWire_61_0_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  vArrayWire_60_0_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vArrayWire_59_0_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  vArrayWire_58_0_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  vArrayWire_57_0_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  vArrayWire_56_0_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  vArrayWire_55_0_r = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  vArrayWire_54_0_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vArrayWire_53_0_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  vArrayWire_52_0_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  vArrayWire_51_0_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  vArrayWire_50_0_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  vArrayWire_49_0_r = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  vArrayWire_48_0_r = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  vArrayWire_47_0_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  vArrayWire_46_0_r = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  vArrayWire_45_0_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  vArrayWire_44_0_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  vArrayWire_43_0_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  vArrayWire_42_0_r = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  vArrayWire_41_0_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  vArrayWire_40_0_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  vArrayWire_39_0_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  vArrayWire_38_0_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vArrayWire_37_0_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  vArrayWire_36_0_r = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  vArrayWire_35_0_r = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  vArrayWire_34_0_r = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  vArrayWire_33_0_r = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  vArrayWire_32_0_r = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  vArrayWire_31_0_r = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  vArrayWire_30_0_r = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  vArrayWire_29_0_r = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  vArrayWire_28_0_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  vArrayWire_27_0_r = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  vArrayWire_26_0_r = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  vArrayWire_25_0_r = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  vArrayWire_24_0_r = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  vArrayWire_23_0_r = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  vArrayWire_22_0_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  vArrayWire_21_0_r = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  vArrayWire_20_0_r = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  vArrayWire_19_0_r = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  vArrayWire_18_0_r = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  vArrayWire_17_0_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  vArrayWire_16_0_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  vArrayWire_15_0_r = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  vArrayWire_14_0_r = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  vArrayWire_13_0_r = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  vArrayWire_12_0_r = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vArrayWire_11_0_r = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  vArrayWire_10_0_r = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  vArrayWire_9_0_r = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  vArrayWire_8_0_r = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  vArrayWire_7_0_r = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  vArrayWire_6_0_r = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  vArrayWire_5_0_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  vArrayWire_4_0_r = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  vArrayWire_3_0_r = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  vArrayWire_2_0_r = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  vArrayWire_1_0_r = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  vArrayWire_0_0_r = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tagArrayWire_63_0_r = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tagArrayWire_62_0_r = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tagArrayWire_61_0_r = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tagArrayWire_60_0_r = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tagArrayWire_59_0_r = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tagArrayWire_58_0_r = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tagArrayWire_57_0_r = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tagArrayWire_56_0_r = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tagArrayWire_55_0_r = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tagArrayWire_54_0_r = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tagArrayWire_53_0_r = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tagArrayWire_52_0_r = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tagArrayWire_51_0_r = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tagArrayWire_50_0_r = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tagArrayWire_49_0_r = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tagArrayWire_48_0_r = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tagArrayWire_47_0_r = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tagArrayWire_46_0_r = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tagArrayWire_45_0_r = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tagArrayWire_44_0_r = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tagArrayWire_43_0_r = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tagArrayWire_42_0_r = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tagArrayWire_41_0_r = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tagArrayWire_40_0_r = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tagArrayWire_39_0_r = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tagArrayWire_38_0_r = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tagArrayWire_37_0_r = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tagArrayWire_36_0_r = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tagArrayWire_35_0_r = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tagArrayWire_34_0_r = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tagArrayWire_33_0_r = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tagArrayWire_32_0_r = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tagArrayWire_31_0_r = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tagArrayWire_30_0_r = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tagArrayWire_29_0_r = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tagArrayWire_28_0_r = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tagArrayWire_27_0_r = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tagArrayWire_26_0_r = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tagArrayWire_25_0_r = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tagArrayWire_24_0_r = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tagArrayWire_23_0_r = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tagArrayWire_22_0_r = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tagArrayWire_21_0_r = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tagArrayWire_20_0_r = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tagArrayWire_19_0_r = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tagArrayWire_18_0_r = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tagArrayWire_17_0_r = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tagArrayWire_16_0_r = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tagArrayWire_15_0_r = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tagArrayWire_14_0_r = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tagArrayWire_13_0_r = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tagArrayWire_12_0_r = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tagArrayWire_11_0_r = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tagArrayWire_10_0_r = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tagArrayWire_9_0_r = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tagArrayWire_8_0_r = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tagArrayWire_7_0_r = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tagArrayWire_6_0_r = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tagArrayWire_5_0_r = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tagArrayWire_4_0_r = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tagArrayWire_3_0_r = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tagArrayWire_2_0_r = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tagArrayWire_1_0_r = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  tagArrayWire_0_0_r = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  vArrayWire_63_1_r = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  vArrayWire_62_1_r = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  vArrayWire_61_1_r = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  vArrayWire_60_1_r = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  vArrayWire_59_1_r = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  vArrayWire_58_1_r = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  vArrayWire_57_1_r = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  vArrayWire_56_1_r = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  vArrayWire_55_1_r = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  vArrayWire_54_1_r = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  vArrayWire_53_1_r = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  vArrayWire_52_1_r = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  vArrayWire_51_1_r = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  vArrayWire_50_1_r = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  vArrayWire_49_1_r = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  vArrayWire_48_1_r = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  vArrayWire_47_1_r = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  vArrayWire_46_1_r = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  vArrayWire_45_1_r = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  vArrayWire_44_1_r = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  vArrayWire_43_1_r = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  vArrayWire_42_1_r = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  vArrayWire_41_1_r = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  vArrayWire_40_1_r = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  vArrayWire_39_1_r = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  vArrayWire_38_1_r = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  vArrayWire_37_1_r = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  vArrayWire_36_1_r = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  vArrayWire_35_1_r = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  vArrayWire_34_1_r = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  vArrayWire_33_1_r = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  vArrayWire_32_1_r = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  vArrayWire_31_1_r = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  vArrayWire_30_1_r = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  vArrayWire_29_1_r = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  vArrayWire_28_1_r = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  vArrayWire_27_1_r = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  vArrayWire_26_1_r = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  vArrayWire_25_1_r = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  vArrayWire_24_1_r = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  vArrayWire_23_1_r = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  vArrayWire_22_1_r = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  vArrayWire_21_1_r = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  vArrayWire_20_1_r = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  vArrayWire_19_1_r = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  vArrayWire_18_1_r = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  vArrayWire_17_1_r = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  vArrayWire_16_1_r = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  vArrayWire_15_1_r = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  vArrayWire_14_1_r = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  vArrayWire_13_1_r = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  vArrayWire_12_1_r = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  vArrayWire_11_1_r = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  vArrayWire_10_1_r = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vArrayWire_9_1_r = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  vArrayWire_8_1_r = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  vArrayWire_7_1_r = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  vArrayWire_6_1_r = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  vArrayWire_5_1_r = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  vArrayWire_4_1_r = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  vArrayWire_3_1_r = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  vArrayWire_2_1_r = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  vArrayWire_1_1_r = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  vArrayWire_0_1_r = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tagArrayWire_63_1_r = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  tagArrayWire_62_1_r = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  tagArrayWire_61_1_r = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  tagArrayWire_60_1_r = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  tagArrayWire_59_1_r = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  tagArrayWire_58_1_r = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  tagArrayWire_57_1_r = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  tagArrayWire_56_1_r = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  tagArrayWire_55_1_r = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  tagArrayWire_54_1_r = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  tagArrayWire_53_1_r = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  tagArrayWire_52_1_r = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  tagArrayWire_51_1_r = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  tagArrayWire_50_1_r = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  tagArrayWire_49_1_r = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  tagArrayWire_48_1_r = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  tagArrayWire_47_1_r = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  tagArrayWire_46_1_r = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  tagArrayWire_45_1_r = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  tagArrayWire_44_1_r = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  tagArrayWire_43_1_r = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  tagArrayWire_42_1_r = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  tagArrayWire_41_1_r = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  tagArrayWire_40_1_r = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  tagArrayWire_39_1_r = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  tagArrayWire_38_1_r = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  tagArrayWire_37_1_r = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  tagArrayWire_36_1_r = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  tagArrayWire_35_1_r = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  tagArrayWire_34_1_r = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  tagArrayWire_33_1_r = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  tagArrayWire_32_1_r = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  tagArrayWire_31_1_r = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  tagArrayWire_30_1_r = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  tagArrayWire_29_1_r = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  tagArrayWire_28_1_r = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  tagArrayWire_27_1_r = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  tagArrayWire_26_1_r = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  tagArrayWire_25_1_r = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  tagArrayWire_24_1_r = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  tagArrayWire_23_1_r = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  tagArrayWire_22_1_r = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  tagArrayWire_21_1_r = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  tagArrayWire_20_1_r = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  tagArrayWire_19_1_r = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  tagArrayWire_18_1_r = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  tagArrayWire_17_1_r = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  tagArrayWire_16_1_r = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  tagArrayWire_15_1_r = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  tagArrayWire_14_1_r = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  tagArrayWire_13_1_r = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  tagArrayWire_12_1_r = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  tagArrayWire_11_1_r = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  tagArrayWire_10_1_r = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  tagArrayWire_9_1_r = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  tagArrayWire_8_1_r = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  tagArrayWire_7_1_r = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  tagArrayWire_6_1_r = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  tagArrayWire_5_1_r = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  tagArrayWire_4_1_r = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  tagArrayWire_3_1_r = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  tagArrayWire_2_1_r = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  tagArrayWire_1_1_r = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  tagArrayWire_0_1_r = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  vArrayWire_63_2_r = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  vArrayWire_62_2_r = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  vArrayWire_61_2_r = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  vArrayWire_60_2_r = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  vArrayWire_59_2_r = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  vArrayWire_58_2_r = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  vArrayWire_57_2_r = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  vArrayWire_56_2_r = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  vArrayWire_55_2_r = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  vArrayWire_54_2_r = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  vArrayWire_53_2_r = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  vArrayWire_52_2_r = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  vArrayWire_51_2_r = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  vArrayWire_50_2_r = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  vArrayWire_49_2_r = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  vArrayWire_48_2_r = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  vArrayWire_47_2_r = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  vArrayWire_46_2_r = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  vArrayWire_45_2_r = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  vArrayWire_44_2_r = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  vArrayWire_43_2_r = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  vArrayWire_42_2_r = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  vArrayWire_41_2_r = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  vArrayWire_40_2_r = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  vArrayWire_39_2_r = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  vArrayWire_38_2_r = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  vArrayWire_37_2_r = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  vArrayWire_36_2_r = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  vArrayWire_35_2_r = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  vArrayWire_34_2_r = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  vArrayWire_33_2_r = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  vArrayWire_32_2_r = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  vArrayWire_31_2_r = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  vArrayWire_30_2_r = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  vArrayWire_29_2_r = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  vArrayWire_28_2_r = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  vArrayWire_27_2_r = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  vArrayWire_26_2_r = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  vArrayWire_25_2_r = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  vArrayWire_24_2_r = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  vArrayWire_23_2_r = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  vArrayWire_22_2_r = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  vArrayWire_21_2_r = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  vArrayWire_20_2_r = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  vArrayWire_19_2_r = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  vArrayWire_18_2_r = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  vArrayWire_17_2_r = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  vArrayWire_16_2_r = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  vArrayWire_15_2_r = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  vArrayWire_14_2_r = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  vArrayWire_13_2_r = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  vArrayWire_12_2_r = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  vArrayWire_11_2_r = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  vArrayWire_10_2_r = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  vArrayWire_9_2_r = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  vArrayWire_8_2_r = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  vArrayWire_7_2_r = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  vArrayWire_6_2_r = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  vArrayWire_5_2_r = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  vArrayWire_4_2_r = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  vArrayWire_3_2_r = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  vArrayWire_2_2_r = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  vArrayWire_1_2_r = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  vArrayWire_0_2_r = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  tagArrayWire_63_2_r = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  tagArrayWire_62_2_r = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  tagArrayWire_61_2_r = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  tagArrayWire_60_2_r = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  tagArrayWire_59_2_r = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  tagArrayWire_58_2_r = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  tagArrayWire_57_2_r = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  tagArrayWire_56_2_r = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  tagArrayWire_55_2_r = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  tagArrayWire_54_2_r = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  tagArrayWire_53_2_r = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  tagArrayWire_52_2_r = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  tagArrayWire_51_2_r = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  tagArrayWire_50_2_r = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  tagArrayWire_49_2_r = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  tagArrayWire_48_2_r = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  tagArrayWire_47_2_r = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  tagArrayWire_46_2_r = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  tagArrayWire_45_2_r = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  tagArrayWire_44_2_r = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  tagArrayWire_43_2_r = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  tagArrayWire_42_2_r = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  tagArrayWire_41_2_r = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  tagArrayWire_40_2_r = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  tagArrayWire_39_2_r = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  tagArrayWire_38_2_r = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  tagArrayWire_37_2_r = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  tagArrayWire_36_2_r = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  tagArrayWire_35_2_r = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  tagArrayWire_34_2_r = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  tagArrayWire_33_2_r = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  tagArrayWire_32_2_r = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  tagArrayWire_31_2_r = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  tagArrayWire_30_2_r = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  tagArrayWire_29_2_r = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  tagArrayWire_28_2_r = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  tagArrayWire_27_2_r = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  tagArrayWire_26_2_r = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  tagArrayWire_25_2_r = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  tagArrayWire_24_2_r = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  tagArrayWire_23_2_r = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  tagArrayWire_22_2_r = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  tagArrayWire_21_2_r = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  tagArrayWire_20_2_r = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  tagArrayWire_19_2_r = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  tagArrayWire_18_2_r = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  tagArrayWire_17_2_r = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  tagArrayWire_16_2_r = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  tagArrayWire_15_2_r = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  tagArrayWire_14_2_r = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  tagArrayWire_13_2_r = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  tagArrayWire_12_2_r = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  tagArrayWire_11_2_r = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  tagArrayWire_10_2_r = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  tagArrayWire_9_2_r = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  tagArrayWire_8_2_r = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  tagArrayWire_7_2_r = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  tagArrayWire_6_2_r = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  tagArrayWire_5_2_r = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  tagArrayWire_4_2_r = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  tagArrayWire_3_2_r = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  tagArrayWire_2_2_r = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  tagArrayWire_1_2_r = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  tagArrayWire_0_2_r = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  vArrayWire_63_3_r = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  vArrayWire_62_3_r = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  vArrayWire_61_3_r = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  vArrayWire_60_3_r = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  vArrayWire_59_3_r = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  vArrayWire_58_3_r = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  vArrayWire_57_3_r = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  vArrayWire_56_3_r = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  vArrayWire_55_3_r = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  vArrayWire_54_3_r = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  vArrayWire_53_3_r = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  vArrayWire_52_3_r = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  vArrayWire_51_3_r = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  vArrayWire_50_3_r = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  vArrayWire_49_3_r = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  vArrayWire_48_3_r = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  vArrayWire_47_3_r = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  vArrayWire_46_3_r = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  vArrayWire_45_3_r = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  vArrayWire_44_3_r = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  vArrayWire_43_3_r = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  vArrayWire_42_3_r = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  vArrayWire_41_3_r = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  vArrayWire_40_3_r = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  vArrayWire_39_3_r = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  vArrayWire_38_3_r = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  vArrayWire_37_3_r = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  vArrayWire_36_3_r = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  vArrayWire_35_3_r = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  vArrayWire_34_3_r = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  vArrayWire_33_3_r = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  vArrayWire_32_3_r = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  vArrayWire_31_3_r = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  vArrayWire_30_3_r = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  vArrayWire_29_3_r = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  vArrayWire_28_3_r = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  vArrayWire_27_3_r = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  vArrayWire_26_3_r = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  vArrayWire_25_3_r = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  vArrayWire_24_3_r = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  vArrayWire_23_3_r = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  vArrayWire_22_3_r = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  vArrayWire_21_3_r = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  vArrayWire_20_3_r = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  vArrayWire_19_3_r = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  vArrayWire_18_3_r = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  vArrayWire_17_3_r = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  vArrayWire_16_3_r = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  vArrayWire_15_3_r = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  vArrayWire_14_3_r = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  vArrayWire_13_3_r = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  vArrayWire_12_3_r = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  vArrayWire_11_3_r = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  vArrayWire_10_3_r = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  vArrayWire_9_3_r = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  vArrayWire_8_3_r = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  vArrayWire_7_3_r = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  vArrayWire_6_3_r = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  vArrayWire_5_3_r = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  vArrayWire_4_3_r = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  vArrayWire_3_3_r = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  vArrayWire_2_3_r = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  vArrayWire_1_3_r = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  vArrayWire_0_3_r = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  tagArrayWire_63_3_r = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  tagArrayWire_62_3_r = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  tagArrayWire_61_3_r = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  tagArrayWire_60_3_r = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  tagArrayWire_59_3_r = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  tagArrayWire_58_3_r = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  tagArrayWire_57_3_r = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  tagArrayWire_56_3_r = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  tagArrayWire_55_3_r = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  tagArrayWire_54_3_r = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  tagArrayWire_53_3_r = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  tagArrayWire_52_3_r = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  tagArrayWire_51_3_r = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  tagArrayWire_50_3_r = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  tagArrayWire_49_3_r = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  tagArrayWire_48_3_r = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  tagArrayWire_47_3_r = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  tagArrayWire_46_3_r = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  tagArrayWire_45_3_r = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  tagArrayWire_44_3_r = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  tagArrayWire_43_3_r = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  tagArrayWire_42_3_r = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  tagArrayWire_41_3_r = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  tagArrayWire_40_3_r = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  tagArrayWire_39_3_r = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  tagArrayWire_38_3_r = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  tagArrayWire_37_3_r = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  tagArrayWire_36_3_r = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  tagArrayWire_35_3_r = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  tagArrayWire_34_3_r = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  tagArrayWire_33_3_r = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  tagArrayWire_32_3_r = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  tagArrayWire_31_3_r = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  tagArrayWire_30_3_r = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  tagArrayWire_29_3_r = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  tagArrayWire_28_3_r = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  tagArrayWire_27_3_r = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  tagArrayWire_26_3_r = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  tagArrayWire_25_3_r = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  tagArrayWire_24_3_r = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  tagArrayWire_23_3_r = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  tagArrayWire_22_3_r = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  tagArrayWire_21_3_r = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  tagArrayWire_20_3_r = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  tagArrayWire_19_3_r = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  tagArrayWire_18_3_r = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  tagArrayWire_17_3_r = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  tagArrayWire_16_3_r = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  tagArrayWire_15_3_r = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  tagArrayWire_14_3_r = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  tagArrayWire_13_3_r = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  tagArrayWire_12_3_r = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  tagArrayWire_11_3_r = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  tagArrayWire_10_3_r = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  tagArrayWire_9_3_r = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  tagArrayWire_8_3_r = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  tagArrayWire_7_3_r = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  tagArrayWire_6_3_r = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  tagArrayWire_5_3_r = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  tagArrayWire_4_3_r = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  tagArrayWire_3_3_r = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  tagArrayWire_2_3_r = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  tagArrayWire_1_3_r = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  tagArrayWire_0_3_r = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  selArrayWire_1_r = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  selArrayWire_0_r = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  selArrayWire_2_r = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  selArrayWire_3_r = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  selArrayWire_4_r = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  selArrayWire_5_r = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  selArrayWire_6_r = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  selArrayWire_7_r = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  selArrayWire_8_r = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  selArrayWire_9_r = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  selArrayWire_10_r = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  selArrayWire_11_r = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  selArrayWire_12_r = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  selArrayWire_13_r = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  selArrayWire_14_r = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  selArrayWire_15_r = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  selArrayWire_16_r = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  selArrayWire_17_r = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  selArrayWire_18_r = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  selArrayWire_19_r = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  selArrayWire_20_r = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  selArrayWire_21_r = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  selArrayWire_22_r = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  selArrayWire_23_r = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  selArrayWire_24_r = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  selArrayWire_25_r = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  selArrayWire_26_r = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  selArrayWire_27_r = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  selArrayWire_28_r = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  selArrayWire_29_r = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  selArrayWire_30_r = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  selArrayWire_31_r = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  selArrayWire_32_r = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  selArrayWire_33_r = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  selArrayWire_34_r = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  selArrayWire_35_r = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  selArrayWire_36_r = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  selArrayWire_37_r = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  selArrayWire_38_r = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  selArrayWire_39_r = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  selArrayWire_40_r = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  selArrayWire_41_r = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  selArrayWire_42_r = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  selArrayWire_43_r = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  selArrayWire_44_r = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  selArrayWire_45_r = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  selArrayWire_46_r = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  selArrayWire_47_r = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  selArrayWire_48_r = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  selArrayWire_49_r = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  selArrayWire_50_r = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  selArrayWire_51_r = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  selArrayWire_52_r = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  selArrayWire_53_r = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  selArrayWire_54_r = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  selArrayWire_55_r = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  selArrayWire_56_r = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  selArrayWire_57_r = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  selArrayWire_58_r = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  selArrayWire_59_r = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  selArrayWire_60_r = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  selArrayWire_61_r = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  selArrayWire_62_r = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  selArrayWire_63_r = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXICache(
  input         clock,
  input         reset,
  input         io_axiIO_awready,
  output        io_axiIO_awvalid,
  output [31:0] io_axiIO_awaddr,
  output [2:0]  io_axiIO_awsize,
  input         io_axiIO_wready,
  output        io_axiIO_wvalid,
  output [63:0] io_axiIO_wdata,
  output [7:0]  io_axiIO_wstrb,
  output        io_axiIO_wlast,
  output        io_axiIO_bready,
  input         io_axiIO_bvalid,
  input         io_axiIO_arready,
  output        io_axiIO_arvalid,
  output [31:0] io_axiIO_araddr,
  output [7:0]  io_axiIO_arlen,
  output [2:0]  io_axiIO_arsize,
  output [1:0]  io_axiIO_arburst,
  output        io_axiIO_rready,
  input         io_axiIO_rvalid,
  input  [63:0] io_axiIO_rdata,
  input         io_axiIO_rlast,
  input         io_cache_ar_valid_o,
  input  [31:0] io_cache_ar_addr_o,
  input  [7:0]  io_cache_ar_len_o,
  output        io_cache_r_valid_i,
  output [63:0] io_cache_r_data_i,
  output        io_cache_r_last_i,
  input         io_cache_w_valid_o,
  output        io_cache_w_ready_i,
  input  [63:0] io_cache_w_data_o,
  input  [31:0] io_cache_w_addr_o,
  input  [7:0]  io_cache_w_mask_o,
  input  [1:0]  io_cache_wsize
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rd_state; // @[AXICache.scala 25:25]
  wire [1:0] r_idle_st = io_cache_ar_valid_o ? 2'h1 : 2'h0; // @[AXICache.scala 26:22]
  wire  _r_req_st_T = io_axiIO_rlast & io_axiIO_rvalid; // @[AXICache.scala 30:22]
  wire [1:0] _r_req_st_T_1 = _r_req_st_T ? 2'h0 : 2'h2; // @[AXICache.scala 29:8]
  wire  isReq = rd_state == 2'h1; // @[AXICache.scala 46:24]
  wire  isData = rd_state == 2'h2; // @[AXICache.scala 47:25]
  wire [1:0] _io_axiIO_arsize_T = isReq ? 2'h3 : 2'h0; // @[AXICache.scala 62:25]
  wire [1:0] valid_c = {io_axiIO_awready,io_axiIO_wready}; // @[Cat.scala 30:58]
  reg [1:0] w_state; // @[AXICache.scala 75:24]
  wire [1:0] w_idle_st = io_cache_w_valid_o ? 2'h1 : 2'h0; // @[AXICache.scala 76:22]
  wire [1:0] _w_req_st_T_1 = 2'h2 == valid_c ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [1:0] w_req_st = 2'h3 == valid_c ? 2'h3 : _w_req_st_T_1; // @[Mux.scala 80:57]
  wire  isWReq = w_state == 2'h1; // @[AXICache.scala 99:24]
  wire  isWData = w_state == 2'h2; // @[AXICache.scala 100:25]
  wire  isWB = w_state == 2'h3; // @[AXICache.scala 101:22]
  wire  _io_axiIO_wvalid_T = isWReq | isWData; // @[AXICache.scala 126:29]
  assign io_axiIO_awvalid = w_state == 2'h1; // @[AXICache.scala 99:24]
  assign io_axiIO_awaddr = isWReq ? io_cache_w_addr_o : 32'h0; // @[AXICache.scala 118:25]
  assign io_axiIO_awsize = {{1'd0}, io_cache_wsize}; // @[AXICache.scala 121:19]
  assign io_axiIO_wvalid = isWReq | isWData; // @[AXICache.scala 126:29]
  assign io_axiIO_wdata = _io_axiIO_wvalid_T ? io_cache_w_data_o : 64'h0; // @[AXICache.scala 127:24]
  assign io_axiIO_wstrb = _io_axiIO_wvalid_T ? io_cache_w_mask_o : 8'h0; // @[AXICache.scala 128:24]
  assign io_axiIO_wlast = isWReq | isWData; // @[AXICache.scala 129:27]
  assign io_axiIO_bready = w_state == 2'h3; // @[AXICache.scala 101:22]
  assign io_axiIO_arvalid = rd_state == 2'h1; // @[AXICache.scala 46:24]
  assign io_axiIO_araddr = isReq ? io_cache_ar_addr_o : 32'h0; // @[AXICache.scala 59:25]
  assign io_axiIO_arlen = isReq ? io_cache_ar_len_o : 8'h0; // @[AXICache.scala 61:23]
  assign io_axiIO_arsize = {{1'd0}, _io_axiIO_arsize_T}; // @[AXICache.scala 62:25]
  assign io_axiIO_arburst = isReq ? 2'h1 : 2'h0; // @[AXICache.scala 63:26]
  assign io_axiIO_rready = isData | isReq; // @[AXICache.scala 66:29]
  assign io_cache_r_valid_i = io_axiIO_rvalid; // @[AXICache.scala 51:22]
  assign io_cache_r_data_i = io_axiIO_rdata; // @[AXICache.scala 52:21]
  assign io_cache_r_last_i = io_axiIO_rlast; // @[AXICache.scala 50:21]
  assign io_cache_w_ready_i = io_axiIO_bvalid & isWB; // @[AXICache.scala 103:41]
  always @(posedge clock) begin
    if (reset) begin // @[AXICache.scala 25:25]
      rd_state <= 2'h0; // @[AXICache.scala 25:25]
    end else if (2'h2 == rd_state) begin // @[Mux.scala 80:57]
      rd_state <= _r_req_st_T_1;
    end else if (2'h1 == rd_state) begin // @[Mux.scala 80:57]
      if (io_axiIO_arready) begin // @[AXICache.scala 27:21]
        rd_state <= _r_req_st_T_1;
      end else begin
        rd_state <= 2'h1;
      end
    end else if (2'h0 == rd_state) begin // @[Mux.scala 80:57]
      rd_state <= r_idle_st;
    end
    if (reset) begin // @[AXICache.scala 75:24]
      w_state <= 2'h0; // @[AXICache.scala 75:24]
    end else if (2'h3 == w_state) begin // @[Mux.scala 80:57]
      if (io_axiIO_bvalid) begin // @[AXICache.scala 86:19]
        w_state <= 2'h0;
      end else begin
        w_state <= 2'h3;
      end
    end else if (2'h2 == w_state) begin // @[Mux.scala 80:57]
      if (io_axiIO_wready) begin // @[AXICache.scala 85:22]
        w_state <= 2'h3;
      end else begin
        w_state <= 2'h2;
      end
    end else if (2'h1 == w_state) begin // @[Mux.scala 80:57]
      w_state <= w_req_st;
    end else begin
      w_state <= w_idle_st;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module arbCpu2DCache(
  input         io_arbIn_valid,
  output        io_arbIn_ready,
  output [63:0] io_arbIn_data_read,
  input  [63:0] io_arbIn_data_write,
  input         io_arbIn_wen,
  input  [31:0] io_arbIn_addr,
  input  [1:0]  io_arbIn_rsize,
  input  [7:0]  io_arbIn_mask,
  output        io_arbMMIO_valid,
  input         io_arbMMIO_ready,
  input  [63:0] io_arbMMIO_data_read,
  output [63:0] io_arbMMIO_data_write,
  output        io_arbMMIO_wen,
  output [31:0] io_arbMMIO_addr,
  output [1:0]  io_arbMMIO_rsize,
  output [7:0]  io_arbMMIO_mask,
  output        io_arbClint_valid,
  input  [63:0] io_arbClint_data_read,
  output [63:0] io_arbClint_data_write,
  output        io_arbClint_wen,
  output [31:0] io_arbClint_addr,
  output        io_arbDCache_valid,
  input         io_arbDCache_ready,
  input  [63:0] io_arbDCache_data_read,
  output [63:0] io_arbDCache_data_write,
  output        io_arbDCache_wen,
  output [31:0] io_arbDCache_addr,
  output [1:0]  io_arbDCache_rsize,
  output [7:0]  io_arbDCache_mask
);
  wire  clinitV = io_arbIn_addr >= 32'h2000000 & io_arbIn_addr < 32'h200bfff; // @[arbCpu2Cache.scala 42:45]
  wire  dCacheV = io_arbIn_addr >= 32'h80000000 & io_arbIn_addr < 32'h8fffffff; // @[arbCpu2Cache.scala 43:44]
  wire  _io_arbMMIO_valid_T_2 = ~clinitV & ~dCacheV; // @[arbCpu2Cache.scala 47:32]
  wire [63:0] _io_arbIn_data_read_T = clinitV ? io_arbClint_data_read : io_arbMMIO_data_read; // @[arbCpu2Cache.scala 57:63]
  assign io_arbIn_ready = clinitV | dCacheV & io_arbDCache_ready | _io_arbMMIO_valid_T_2 & io_arbMMIO_ready; // @[arbCpu2Cache.scala 56:86]
  assign io_arbIn_data_read = dCacheV ? io_arbDCache_data_read : _io_arbIn_data_read_T; // @[arbCpu2Cache.scala 57:27]
  assign io_arbMMIO_valid = ~clinitV & ~dCacheV & io_arbIn_valid; // @[arbCpu2Cache.scala 47:44]
  assign io_arbMMIO_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 50:23]
  assign io_arbMMIO_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 50:23]
  assign io_arbClint_valid = clinitV & io_arbIn_valid; // @[arbCpu2Cache.scala 45:32]
  assign io_arbClint_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 51:24]
  assign io_arbClint_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 51:24]
  assign io_arbClint_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 51:24]
  assign io_arbDCache_valid = dCacheV & io_arbIn_valid; // @[arbCpu2Cache.scala 46:33]
  assign io_arbDCache_data_write = io_arbIn_data_write; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_wen = io_arbIn_wen; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_addr = io_arbIn_addr; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_rsize = io_arbIn_rsize; // @[arbCpu2Cache.scala 52:25]
  assign io_arbDCache_mask = io_arbIn_mask; // @[arbCpu2Cache.scala 52:25]
endmodule
module mmioCache(
  input         clock,
  input         reset,
  input         io_block,
  input         io_mmioIn_valid,
  output        io_mmioIn_ready,
  output [63:0] io_mmioIn_data_read,
  input  [63:0] io_mmioIn_data_write,
  input         io_mmioIn_wen,
  input  [31:0] io_mmioIn_addr,
  input  [1:0]  io_mmioIn_rsize,
  input  [7:0]  io_mmioIn_mask,
  output        io_mmioOut_valid,
  input         io_mmioOut_ready,
  input  [63:0] io_mmioOut_data_read,
  output [63:0] io_mmioOut_data_write,
  output        io_mmioOut_wen,
  output [31:0] io_mmioOut_addr,
  output [1:0]  io_mmioOut_rsize,
  output [7:0]  io_mmioOut_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] idleMux = io_mmioIn_valid ? 2'h1 : 2'h0; // @[mmioCache.scala 14:20]
  reg [1:0] state; // @[mmioCache.scala 17:22]
  wire  isIdle = state == 2'h0; // @[mmioCache.scala 27:22]
  reg [63:0] io_mmioIn_data_read_r; // @[Reg.scala 27:20]
  assign io_mmioIn_ready = state == 2'h2; // @[mmioCache.scala 29:22]
  assign io_mmioIn_data_read = io_mmioIn_data_read_r; // @[mmioCache.scala 38:23]
  assign io_mmioOut_valid = isIdle & io_mmioIn_valid; // @[mmioCache.scala 31:30]
  assign io_mmioOut_data_write = io_mmioIn_data_write; // @[mmioCache.scala 35:25]
  assign io_mmioOut_wen = io_mmioIn_wen; // @[mmioCache.scala 32:18]
  assign io_mmioOut_addr = io_mmioIn_addr; // @[mmioCache.scala 33:19]
  assign io_mmioOut_rsize = io_mmioIn_rsize; // @[mmioCache.scala 36:20]
  assign io_mmioOut_mask = io_mmioIn_mask; // @[mmioCache.scala 34:19]
  always @(posedge clock) begin
    if (reset) begin // @[mmioCache.scala 17:22]
      state <= 2'h0; // @[mmioCache.scala 17:22]
    end else if (2'h2 == state) begin // @[Mux.scala 80:57]
      if (io_block) begin // @[mmioCache.scala 16:20]
        state <= 2'h2;
      end else begin
        state <= 2'h0;
      end
    end else if (2'h1 == state) begin // @[Mux.scala 80:57]
      if (io_mmioOut_ready) begin // @[mmioCache.scala 15:20]
        state <= 2'h2;
      end else begin
        state <= 2'h1;
      end
    end else if (2'h0 == state) begin // @[Mux.scala 80:57]
      state <= idleMux;
    end else begin
      state <= 2'h0;
    end
    if (reset) begin // @[Reg.scala 27:20]
      io_mmioIn_data_read_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (io_mmioOut_ready) begin // @[Reg.scala 28:19]
      io_mmioIn_data_read_r <= io_mmioOut_data_read; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  io_mmioIn_data_read_r = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Dcache(
  input          clock,
  input          reset,
  output         io_cacheOut_ar_valid_o,
  output [31:0]  io_cacheOut_ar_addr_o,
  output [7:0]   io_cacheOut_ar_len_o,
  input          io_cacheOut_r_valid_i,
  input  [63:0]  io_cacheOut_r_data_i,
  input          io_cacheOut_r_last_i,
  output         io_cacheOut_w_valid_o,
  input          io_cacheOut_w_ready_i,
  output [63:0]  io_cacheOut_w_data_o,
  output [31:0]  io_cacheOut_w_addr_o,
  output [7:0]   io_cacheOut_w_mask_o,
  output [1:0]   io_cacheOut_wsize,
  input          io_cacheIn_valid,
  output         io_cacheIn_ready,
  output [63:0]  io_cacheIn_data_read,
  input  [63:0]  io_cacheIn_data_write,
  input          io_cacheIn_wen,
  input  [31:0]  io_cacheIn_addr,
  input  [1:0]   io_cacheIn_rsize,
  input  [7:0]   io_cacheIn_mask,
  output         io_SRAMIO_0_cen,
  output         io_SRAMIO_0_wen,
  output [127:0] io_SRAMIO_0_wdata,
  output [5:0]   io_SRAMIO_0_addr,
  output [127:0] io_SRAMIO_0_wmask,
  input  [127:0] io_SRAMIO_0_rdata,
  output         io_SRAMIO_1_cen,
  output         io_SRAMIO_1_wen,
  output [127:0] io_SRAMIO_1_wdata,
  output [5:0]   io_SRAMIO_1_addr,
  output [127:0] io_SRAMIO_1_wmask,
  input  [127:0] io_SRAMIO_1_rdata,
  output         io_SRAMIO_2_cen,
  output         io_SRAMIO_2_wen,
  output [127:0] io_SRAMIO_2_wdata,
  output [5:0]   io_SRAMIO_2_addr,
  output [127:0] io_SRAMIO_2_wmask,
  input  [127:0] io_SRAMIO_2_rdata,
  output         io_SRAMIO_3_cen,
  output         io_SRAMIO_3_wen,
  output [127:0] io_SRAMIO_3_wdata,
  output [5:0]   io_SRAMIO_3_addr,
  output [127:0] io_SRAMIO_3_wmask,
  input  [127:0] io_SRAMIO_3_rdata,
  input          io_block
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] offset = io_cacheIn_addr[3:0]; // @[Cache.scala 173:31]
  wire [5:0] index = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  wire [21:0] tag = io_cacheIn_addr[31:10]; // @[Cache.scala 175:28]
  reg [1:0] cacheState; // @[Cache.scala 178:27]
  wire  _IdleMux_T_1 = io_cacheIn_valid & ~io_block; // @[Cache.scala 182:22]
  wire  _vMuxOut_T_124 = 6'h3f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_63_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_122 = 6'h3e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_62_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_120 = 6'h3d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_61_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_118 = 6'h3c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_60_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_116 = 6'h3b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_59_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_114 = 6'h3a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_58_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_112 = 6'h39 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_57_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_110 = 6'h38 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_56_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_108 = 6'h37 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_55_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_106 = 6'h36 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_54_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_104 = 6'h35 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_53_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_102 = 6'h34 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_52_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_100 = 6'h33 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_51_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_98 = 6'h32 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_50_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_96 = 6'h31 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_49_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_94 = 6'h30 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_48_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_92 = 6'h2f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_47_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_90 = 6'h2e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_46_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_88 = 6'h2d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_45_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_86 = 6'h2c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_44_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_84 = 6'h2b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_43_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_82 = 6'h2a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_42_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_80 = 6'h29 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_41_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_78 = 6'h28 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_40_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_76 = 6'h27 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_39_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_74 = 6'h26 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_38_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_72 = 6'h25 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_37_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_70 = 6'h24 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_36_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_68 = 6'h23 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_35_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_66 = 6'h22 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_34_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_64 = 6'h21 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_33_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_62 = 6'h20 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_32_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_60 = 6'h1f == index; // @[Mux.scala 80:60]
  reg  vArrayWire_31_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_58 = 6'h1e == index; // @[Mux.scala 80:60]
  reg  vArrayWire_30_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_56 = 6'h1d == index; // @[Mux.scala 80:60]
  reg  vArrayWire_29_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_54 = 6'h1c == index; // @[Mux.scala 80:60]
  reg  vArrayWire_28_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_52 = 6'h1b == index; // @[Mux.scala 80:60]
  reg  vArrayWire_27_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_50 = 6'h1a == index; // @[Mux.scala 80:60]
  reg  vArrayWire_26_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_48 = 6'h19 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_25_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_46 = 6'h18 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_24_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_44 = 6'h17 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_23_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_42 = 6'h16 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_22_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_40 = 6'h15 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_21_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_38 = 6'h14 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_20_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_36 = 6'h13 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_19_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_34 = 6'h12 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_18_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_32 = 6'h11 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_17_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_30 = 6'h10 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_16_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_28 = 6'hf == index; // @[Mux.scala 80:60]
  reg  vArrayWire_15_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_26 = 6'he == index; // @[Mux.scala 80:60]
  reg  vArrayWire_14_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_24 = 6'hd == index; // @[Mux.scala 80:60]
  reg  vArrayWire_13_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_22 = 6'hc == index; // @[Mux.scala 80:60]
  reg  vArrayWire_12_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_20 = 6'hb == index; // @[Mux.scala 80:60]
  reg  vArrayWire_11_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_18 = 6'ha == index; // @[Mux.scala 80:60]
  reg  vArrayWire_10_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_16 = 6'h9 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_9_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_14 = 6'h8 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_8_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_12 = 6'h7 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_7_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_10 = 6'h6 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_6_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_8 = 6'h5 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_5_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_6 = 6'h4 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_4_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_4 = 6'h3 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_3_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_2 = 6'h2 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_2_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T = 6'h1 == index; // @[Mux.scala 80:60]
  reg  vArrayWire_1_0_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_0_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_0 = 6'h1 == index ? vArrayWire_1_0_r : vArrayWire_0_0_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_0 = 6'h2 == index ? vArrayWire_2_0_r : _vMuxOut_T_1_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_0 = 6'h3 == index ? vArrayWire_3_0_r : _vMuxOut_T_3_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_0 = 6'h4 == index ? vArrayWire_4_0_r : _vMuxOut_T_5_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_0 = 6'h5 == index ? vArrayWire_5_0_r : _vMuxOut_T_7_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_0 = 6'h6 == index ? vArrayWire_6_0_r : _vMuxOut_T_9_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_0 = 6'h7 == index ? vArrayWire_7_0_r : _vMuxOut_T_11_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_0 = 6'h8 == index ? vArrayWire_8_0_r : _vMuxOut_T_13_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_0 = 6'h9 == index ? vArrayWire_9_0_r : _vMuxOut_T_15_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_0 = 6'ha == index ? vArrayWire_10_0_r : _vMuxOut_T_17_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_0 = 6'hb == index ? vArrayWire_11_0_r : _vMuxOut_T_19_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_0 = 6'hc == index ? vArrayWire_12_0_r : _vMuxOut_T_21_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_0 = 6'hd == index ? vArrayWire_13_0_r : _vMuxOut_T_23_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_0 = 6'he == index ? vArrayWire_14_0_r : _vMuxOut_T_25_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_0 = 6'hf == index ? vArrayWire_15_0_r : _vMuxOut_T_27_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_0 = 6'h10 == index ? vArrayWire_16_0_r : _vMuxOut_T_29_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_0 = 6'h11 == index ? vArrayWire_17_0_r : _vMuxOut_T_31_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_0 = 6'h12 == index ? vArrayWire_18_0_r : _vMuxOut_T_33_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_0 = 6'h13 == index ? vArrayWire_19_0_r : _vMuxOut_T_35_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_0 = 6'h14 == index ? vArrayWire_20_0_r : _vMuxOut_T_37_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_0 = 6'h15 == index ? vArrayWire_21_0_r : _vMuxOut_T_39_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_0 = 6'h16 == index ? vArrayWire_22_0_r : _vMuxOut_T_41_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_0 = 6'h17 == index ? vArrayWire_23_0_r : _vMuxOut_T_43_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_0 = 6'h18 == index ? vArrayWire_24_0_r : _vMuxOut_T_45_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_0 = 6'h19 == index ? vArrayWire_25_0_r : _vMuxOut_T_47_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_0 = 6'h1a == index ? vArrayWire_26_0_r : _vMuxOut_T_49_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_0 = 6'h1b == index ? vArrayWire_27_0_r : _vMuxOut_T_51_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_0 = 6'h1c == index ? vArrayWire_28_0_r : _vMuxOut_T_53_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_0 = 6'h1d == index ? vArrayWire_29_0_r : _vMuxOut_T_55_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_0 = 6'h1e == index ? vArrayWire_30_0_r : _vMuxOut_T_57_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_0 = 6'h1f == index ? vArrayWire_31_0_r : _vMuxOut_T_59_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_0 = 6'h20 == index ? vArrayWire_32_0_r : _vMuxOut_T_61_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_0 = 6'h21 == index ? vArrayWire_33_0_r : _vMuxOut_T_63_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_0 = 6'h22 == index ? vArrayWire_34_0_r : _vMuxOut_T_65_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_0 = 6'h23 == index ? vArrayWire_35_0_r : _vMuxOut_T_67_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_0 = 6'h24 == index ? vArrayWire_36_0_r : _vMuxOut_T_69_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_0 = 6'h25 == index ? vArrayWire_37_0_r : _vMuxOut_T_71_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_0 = 6'h26 == index ? vArrayWire_38_0_r : _vMuxOut_T_73_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_0 = 6'h27 == index ? vArrayWire_39_0_r : _vMuxOut_T_75_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_0 = 6'h28 == index ? vArrayWire_40_0_r : _vMuxOut_T_77_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_0 = 6'h29 == index ? vArrayWire_41_0_r : _vMuxOut_T_79_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_0 = 6'h2a == index ? vArrayWire_42_0_r : _vMuxOut_T_81_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_0 = 6'h2b == index ? vArrayWire_43_0_r : _vMuxOut_T_83_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_0 = 6'h2c == index ? vArrayWire_44_0_r : _vMuxOut_T_85_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_0 = 6'h2d == index ? vArrayWire_45_0_r : _vMuxOut_T_87_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_0 = 6'h2e == index ? vArrayWire_46_0_r : _vMuxOut_T_89_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_0 = 6'h2f == index ? vArrayWire_47_0_r : _vMuxOut_T_91_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_0 = 6'h30 == index ? vArrayWire_48_0_r : _vMuxOut_T_93_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_0 = 6'h31 == index ? vArrayWire_49_0_r : _vMuxOut_T_95_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_0 = 6'h32 == index ? vArrayWire_50_0_r : _vMuxOut_T_97_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_0 = 6'h33 == index ? vArrayWire_51_0_r : _vMuxOut_T_99_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_0 = 6'h34 == index ? vArrayWire_52_0_r : _vMuxOut_T_101_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_0 = 6'h35 == index ? vArrayWire_53_0_r : _vMuxOut_T_103_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_0 = 6'h36 == index ? vArrayWire_54_0_r : _vMuxOut_T_105_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_0 = 6'h37 == index ? vArrayWire_55_0_r : _vMuxOut_T_107_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_0 = 6'h38 == index ? vArrayWire_56_0_r : _vMuxOut_T_109_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_0 = 6'h39 == index ? vArrayWire_57_0_r : _vMuxOut_T_111_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_0 = 6'h3a == index ? vArrayWire_58_0_r : _vMuxOut_T_113_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_0 = 6'h3b == index ? vArrayWire_59_0_r : _vMuxOut_T_115_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_0 = 6'h3c == index ? vArrayWire_60_0_r : _vMuxOut_T_117_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_0 = 6'h3d == index ? vArrayWire_61_0_r : _vMuxOut_T_119_0; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_0 = 6'h3e == index ? vArrayWire_62_0_r : _vMuxOut_T_121_0; // @[Mux.scala 80:57]
  wire  vMuxOut_0 = 6'h3f == index ? vArrayWire_63_0_r : _vMuxOut_T_123_0; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_0_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_0_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_0 = 6'h1 == index ? tagArrayWire_1_0_r : tagArrayWire_0_0_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_0 = 6'h2 == index ? tagArrayWire_2_0_r : _tagMuxOut_T_1_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_0 = 6'h3 == index ? tagArrayWire_3_0_r : _tagMuxOut_T_3_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_0 = 6'h4 == index ? tagArrayWire_4_0_r : _tagMuxOut_T_5_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_0 = 6'h5 == index ? tagArrayWire_5_0_r : _tagMuxOut_T_7_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_0 = 6'h6 == index ? tagArrayWire_6_0_r : _tagMuxOut_T_9_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_0 = 6'h7 == index ? tagArrayWire_7_0_r : _tagMuxOut_T_11_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_0 = 6'h8 == index ? tagArrayWire_8_0_r : _tagMuxOut_T_13_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_0 = 6'h9 == index ? tagArrayWire_9_0_r : _tagMuxOut_T_15_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_0 = 6'ha == index ? tagArrayWire_10_0_r : _tagMuxOut_T_17_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_0 = 6'hb == index ? tagArrayWire_11_0_r : _tagMuxOut_T_19_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_0 = 6'hc == index ? tagArrayWire_12_0_r : _tagMuxOut_T_21_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_0 = 6'hd == index ? tagArrayWire_13_0_r : _tagMuxOut_T_23_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_0 = 6'he == index ? tagArrayWire_14_0_r : _tagMuxOut_T_25_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_0 = 6'hf == index ? tagArrayWire_15_0_r : _tagMuxOut_T_27_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_0 = 6'h10 == index ? tagArrayWire_16_0_r : _tagMuxOut_T_29_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_0 = 6'h11 == index ? tagArrayWire_17_0_r : _tagMuxOut_T_31_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_0 = 6'h12 == index ? tagArrayWire_18_0_r : _tagMuxOut_T_33_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_0 = 6'h13 == index ? tagArrayWire_19_0_r : _tagMuxOut_T_35_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_0 = 6'h14 == index ? tagArrayWire_20_0_r : _tagMuxOut_T_37_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_0 = 6'h15 == index ? tagArrayWire_21_0_r : _tagMuxOut_T_39_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_0 = 6'h16 == index ? tagArrayWire_22_0_r : _tagMuxOut_T_41_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_0 = 6'h17 == index ? tagArrayWire_23_0_r : _tagMuxOut_T_43_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_0 = 6'h18 == index ? tagArrayWire_24_0_r : _tagMuxOut_T_45_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_0 = 6'h19 == index ? tagArrayWire_25_0_r : _tagMuxOut_T_47_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_0 = 6'h1a == index ? tagArrayWire_26_0_r : _tagMuxOut_T_49_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_0 = 6'h1b == index ? tagArrayWire_27_0_r : _tagMuxOut_T_51_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_0 = 6'h1c == index ? tagArrayWire_28_0_r : _tagMuxOut_T_53_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_0 = 6'h1d == index ? tagArrayWire_29_0_r : _tagMuxOut_T_55_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_0 = 6'h1e == index ? tagArrayWire_30_0_r : _tagMuxOut_T_57_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_0 = 6'h1f == index ? tagArrayWire_31_0_r : _tagMuxOut_T_59_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_0 = 6'h20 == index ? tagArrayWire_32_0_r : _tagMuxOut_T_61_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_0 = 6'h21 == index ? tagArrayWire_33_0_r : _tagMuxOut_T_63_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_0 = 6'h22 == index ? tagArrayWire_34_0_r : _tagMuxOut_T_65_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_0 = 6'h23 == index ? tagArrayWire_35_0_r : _tagMuxOut_T_67_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_0 = 6'h24 == index ? tagArrayWire_36_0_r : _tagMuxOut_T_69_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_0 = 6'h25 == index ? tagArrayWire_37_0_r : _tagMuxOut_T_71_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_0 = 6'h26 == index ? tagArrayWire_38_0_r : _tagMuxOut_T_73_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_0 = 6'h27 == index ? tagArrayWire_39_0_r : _tagMuxOut_T_75_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_0 = 6'h28 == index ? tagArrayWire_40_0_r : _tagMuxOut_T_77_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_0 = 6'h29 == index ? tagArrayWire_41_0_r : _tagMuxOut_T_79_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_0 = 6'h2a == index ? tagArrayWire_42_0_r : _tagMuxOut_T_81_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_0 = 6'h2b == index ? tagArrayWire_43_0_r : _tagMuxOut_T_83_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_0 = 6'h2c == index ? tagArrayWire_44_0_r : _tagMuxOut_T_85_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_0 = 6'h2d == index ? tagArrayWire_45_0_r : _tagMuxOut_T_87_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_0 = 6'h2e == index ? tagArrayWire_46_0_r : _tagMuxOut_T_89_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_0 = 6'h2f == index ? tagArrayWire_47_0_r : _tagMuxOut_T_91_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_0 = 6'h30 == index ? tagArrayWire_48_0_r : _tagMuxOut_T_93_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_0 = 6'h31 == index ? tagArrayWire_49_0_r : _tagMuxOut_T_95_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_0 = 6'h32 == index ? tagArrayWire_50_0_r : _tagMuxOut_T_97_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_0 = 6'h33 == index ? tagArrayWire_51_0_r : _tagMuxOut_T_99_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_0 = 6'h34 == index ? tagArrayWire_52_0_r : _tagMuxOut_T_101_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_0 = 6'h35 == index ? tagArrayWire_53_0_r : _tagMuxOut_T_103_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_0 = 6'h36 == index ? tagArrayWire_54_0_r : _tagMuxOut_T_105_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_0 = 6'h37 == index ? tagArrayWire_55_0_r : _tagMuxOut_T_107_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_0 = 6'h38 == index ? tagArrayWire_56_0_r : _tagMuxOut_T_109_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_0 = 6'h39 == index ? tagArrayWire_57_0_r : _tagMuxOut_T_111_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_0 = 6'h3a == index ? tagArrayWire_58_0_r : _tagMuxOut_T_113_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_0 = 6'h3b == index ? tagArrayWire_59_0_r : _tagMuxOut_T_115_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_0 = 6'h3c == index ? tagArrayWire_60_0_r : _tagMuxOut_T_117_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_0 = 6'h3d == index ? tagArrayWire_61_0_r : _tagMuxOut_T_119_0; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_0 = 6'h3e == index ? tagArrayWire_62_0_r : _tagMuxOut_T_121_0; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_0 = 6'h3f == index ? tagArrayWire_63_0_r : _tagMuxOut_T_123_0; // @[Mux.scala 80:57]
  wire  hitArray_0 = vMuxOut_0 & tagMuxOut_0 == tag; // @[Cache.scala 243:60]
  reg  vArrayWire_63_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_1_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_1_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_1 = 6'h1 == index ? vArrayWire_1_1_r : vArrayWire_0_1_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_1 = 6'h2 == index ? vArrayWire_2_1_r : _vMuxOut_T_1_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_1 = 6'h3 == index ? vArrayWire_3_1_r : _vMuxOut_T_3_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_1 = 6'h4 == index ? vArrayWire_4_1_r : _vMuxOut_T_5_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_1 = 6'h5 == index ? vArrayWire_5_1_r : _vMuxOut_T_7_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_1 = 6'h6 == index ? vArrayWire_6_1_r : _vMuxOut_T_9_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_1 = 6'h7 == index ? vArrayWire_7_1_r : _vMuxOut_T_11_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_1 = 6'h8 == index ? vArrayWire_8_1_r : _vMuxOut_T_13_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_1 = 6'h9 == index ? vArrayWire_9_1_r : _vMuxOut_T_15_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_1 = 6'ha == index ? vArrayWire_10_1_r : _vMuxOut_T_17_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_1 = 6'hb == index ? vArrayWire_11_1_r : _vMuxOut_T_19_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_1 = 6'hc == index ? vArrayWire_12_1_r : _vMuxOut_T_21_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_1 = 6'hd == index ? vArrayWire_13_1_r : _vMuxOut_T_23_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_1 = 6'he == index ? vArrayWire_14_1_r : _vMuxOut_T_25_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_1 = 6'hf == index ? vArrayWire_15_1_r : _vMuxOut_T_27_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_1 = 6'h10 == index ? vArrayWire_16_1_r : _vMuxOut_T_29_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_1 = 6'h11 == index ? vArrayWire_17_1_r : _vMuxOut_T_31_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_1 = 6'h12 == index ? vArrayWire_18_1_r : _vMuxOut_T_33_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_1 = 6'h13 == index ? vArrayWire_19_1_r : _vMuxOut_T_35_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_1 = 6'h14 == index ? vArrayWire_20_1_r : _vMuxOut_T_37_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_1 = 6'h15 == index ? vArrayWire_21_1_r : _vMuxOut_T_39_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_1 = 6'h16 == index ? vArrayWire_22_1_r : _vMuxOut_T_41_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_1 = 6'h17 == index ? vArrayWire_23_1_r : _vMuxOut_T_43_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_1 = 6'h18 == index ? vArrayWire_24_1_r : _vMuxOut_T_45_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_1 = 6'h19 == index ? vArrayWire_25_1_r : _vMuxOut_T_47_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_1 = 6'h1a == index ? vArrayWire_26_1_r : _vMuxOut_T_49_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_1 = 6'h1b == index ? vArrayWire_27_1_r : _vMuxOut_T_51_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_1 = 6'h1c == index ? vArrayWire_28_1_r : _vMuxOut_T_53_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_1 = 6'h1d == index ? vArrayWire_29_1_r : _vMuxOut_T_55_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_1 = 6'h1e == index ? vArrayWire_30_1_r : _vMuxOut_T_57_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_1 = 6'h1f == index ? vArrayWire_31_1_r : _vMuxOut_T_59_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_1 = 6'h20 == index ? vArrayWire_32_1_r : _vMuxOut_T_61_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_1 = 6'h21 == index ? vArrayWire_33_1_r : _vMuxOut_T_63_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_1 = 6'h22 == index ? vArrayWire_34_1_r : _vMuxOut_T_65_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_1 = 6'h23 == index ? vArrayWire_35_1_r : _vMuxOut_T_67_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_1 = 6'h24 == index ? vArrayWire_36_1_r : _vMuxOut_T_69_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_1 = 6'h25 == index ? vArrayWire_37_1_r : _vMuxOut_T_71_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_1 = 6'h26 == index ? vArrayWire_38_1_r : _vMuxOut_T_73_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_1 = 6'h27 == index ? vArrayWire_39_1_r : _vMuxOut_T_75_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_1 = 6'h28 == index ? vArrayWire_40_1_r : _vMuxOut_T_77_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_1 = 6'h29 == index ? vArrayWire_41_1_r : _vMuxOut_T_79_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_1 = 6'h2a == index ? vArrayWire_42_1_r : _vMuxOut_T_81_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_1 = 6'h2b == index ? vArrayWire_43_1_r : _vMuxOut_T_83_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_1 = 6'h2c == index ? vArrayWire_44_1_r : _vMuxOut_T_85_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_1 = 6'h2d == index ? vArrayWire_45_1_r : _vMuxOut_T_87_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_1 = 6'h2e == index ? vArrayWire_46_1_r : _vMuxOut_T_89_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_1 = 6'h2f == index ? vArrayWire_47_1_r : _vMuxOut_T_91_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_1 = 6'h30 == index ? vArrayWire_48_1_r : _vMuxOut_T_93_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_1 = 6'h31 == index ? vArrayWire_49_1_r : _vMuxOut_T_95_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_1 = 6'h32 == index ? vArrayWire_50_1_r : _vMuxOut_T_97_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_1 = 6'h33 == index ? vArrayWire_51_1_r : _vMuxOut_T_99_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_1 = 6'h34 == index ? vArrayWire_52_1_r : _vMuxOut_T_101_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_1 = 6'h35 == index ? vArrayWire_53_1_r : _vMuxOut_T_103_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_1 = 6'h36 == index ? vArrayWire_54_1_r : _vMuxOut_T_105_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_1 = 6'h37 == index ? vArrayWire_55_1_r : _vMuxOut_T_107_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_1 = 6'h38 == index ? vArrayWire_56_1_r : _vMuxOut_T_109_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_1 = 6'h39 == index ? vArrayWire_57_1_r : _vMuxOut_T_111_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_1 = 6'h3a == index ? vArrayWire_58_1_r : _vMuxOut_T_113_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_1 = 6'h3b == index ? vArrayWire_59_1_r : _vMuxOut_T_115_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_1 = 6'h3c == index ? vArrayWire_60_1_r : _vMuxOut_T_117_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_1 = 6'h3d == index ? vArrayWire_61_1_r : _vMuxOut_T_119_1; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_1 = 6'h3e == index ? vArrayWire_62_1_r : _vMuxOut_T_121_1; // @[Mux.scala 80:57]
  wire  vMuxOut_1 = 6'h3f == index ? vArrayWire_63_1_r : _vMuxOut_T_123_1; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_1_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_1_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_1 = 6'h1 == index ? tagArrayWire_1_1_r : tagArrayWire_0_1_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_1 = 6'h2 == index ? tagArrayWire_2_1_r : _tagMuxOut_T_1_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_1 = 6'h3 == index ? tagArrayWire_3_1_r : _tagMuxOut_T_3_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_1 = 6'h4 == index ? tagArrayWire_4_1_r : _tagMuxOut_T_5_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_1 = 6'h5 == index ? tagArrayWire_5_1_r : _tagMuxOut_T_7_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_1 = 6'h6 == index ? tagArrayWire_6_1_r : _tagMuxOut_T_9_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_1 = 6'h7 == index ? tagArrayWire_7_1_r : _tagMuxOut_T_11_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_1 = 6'h8 == index ? tagArrayWire_8_1_r : _tagMuxOut_T_13_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_1 = 6'h9 == index ? tagArrayWire_9_1_r : _tagMuxOut_T_15_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_1 = 6'ha == index ? tagArrayWire_10_1_r : _tagMuxOut_T_17_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_1 = 6'hb == index ? tagArrayWire_11_1_r : _tagMuxOut_T_19_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_1 = 6'hc == index ? tagArrayWire_12_1_r : _tagMuxOut_T_21_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_1 = 6'hd == index ? tagArrayWire_13_1_r : _tagMuxOut_T_23_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_1 = 6'he == index ? tagArrayWire_14_1_r : _tagMuxOut_T_25_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_1 = 6'hf == index ? tagArrayWire_15_1_r : _tagMuxOut_T_27_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_1 = 6'h10 == index ? tagArrayWire_16_1_r : _tagMuxOut_T_29_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_1 = 6'h11 == index ? tagArrayWire_17_1_r : _tagMuxOut_T_31_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_1 = 6'h12 == index ? tagArrayWire_18_1_r : _tagMuxOut_T_33_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_1 = 6'h13 == index ? tagArrayWire_19_1_r : _tagMuxOut_T_35_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_1 = 6'h14 == index ? tagArrayWire_20_1_r : _tagMuxOut_T_37_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_1 = 6'h15 == index ? tagArrayWire_21_1_r : _tagMuxOut_T_39_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_1 = 6'h16 == index ? tagArrayWire_22_1_r : _tagMuxOut_T_41_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_1 = 6'h17 == index ? tagArrayWire_23_1_r : _tagMuxOut_T_43_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_1 = 6'h18 == index ? tagArrayWire_24_1_r : _tagMuxOut_T_45_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_1 = 6'h19 == index ? tagArrayWire_25_1_r : _tagMuxOut_T_47_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_1 = 6'h1a == index ? tagArrayWire_26_1_r : _tagMuxOut_T_49_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_1 = 6'h1b == index ? tagArrayWire_27_1_r : _tagMuxOut_T_51_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_1 = 6'h1c == index ? tagArrayWire_28_1_r : _tagMuxOut_T_53_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_1 = 6'h1d == index ? tagArrayWire_29_1_r : _tagMuxOut_T_55_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_1 = 6'h1e == index ? tagArrayWire_30_1_r : _tagMuxOut_T_57_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_1 = 6'h1f == index ? tagArrayWire_31_1_r : _tagMuxOut_T_59_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_1 = 6'h20 == index ? tagArrayWire_32_1_r : _tagMuxOut_T_61_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_1 = 6'h21 == index ? tagArrayWire_33_1_r : _tagMuxOut_T_63_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_1 = 6'h22 == index ? tagArrayWire_34_1_r : _tagMuxOut_T_65_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_1 = 6'h23 == index ? tagArrayWire_35_1_r : _tagMuxOut_T_67_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_1 = 6'h24 == index ? tagArrayWire_36_1_r : _tagMuxOut_T_69_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_1 = 6'h25 == index ? tagArrayWire_37_1_r : _tagMuxOut_T_71_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_1 = 6'h26 == index ? tagArrayWire_38_1_r : _tagMuxOut_T_73_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_1 = 6'h27 == index ? tagArrayWire_39_1_r : _tagMuxOut_T_75_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_1 = 6'h28 == index ? tagArrayWire_40_1_r : _tagMuxOut_T_77_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_1 = 6'h29 == index ? tagArrayWire_41_1_r : _tagMuxOut_T_79_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_1 = 6'h2a == index ? tagArrayWire_42_1_r : _tagMuxOut_T_81_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_1 = 6'h2b == index ? tagArrayWire_43_1_r : _tagMuxOut_T_83_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_1 = 6'h2c == index ? tagArrayWire_44_1_r : _tagMuxOut_T_85_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_1 = 6'h2d == index ? tagArrayWire_45_1_r : _tagMuxOut_T_87_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_1 = 6'h2e == index ? tagArrayWire_46_1_r : _tagMuxOut_T_89_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_1 = 6'h2f == index ? tagArrayWire_47_1_r : _tagMuxOut_T_91_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_1 = 6'h30 == index ? tagArrayWire_48_1_r : _tagMuxOut_T_93_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_1 = 6'h31 == index ? tagArrayWire_49_1_r : _tagMuxOut_T_95_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_1 = 6'h32 == index ? tagArrayWire_50_1_r : _tagMuxOut_T_97_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_1 = 6'h33 == index ? tagArrayWire_51_1_r : _tagMuxOut_T_99_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_1 = 6'h34 == index ? tagArrayWire_52_1_r : _tagMuxOut_T_101_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_1 = 6'h35 == index ? tagArrayWire_53_1_r : _tagMuxOut_T_103_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_1 = 6'h36 == index ? tagArrayWire_54_1_r : _tagMuxOut_T_105_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_1 = 6'h37 == index ? tagArrayWire_55_1_r : _tagMuxOut_T_107_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_1 = 6'h38 == index ? tagArrayWire_56_1_r : _tagMuxOut_T_109_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_1 = 6'h39 == index ? tagArrayWire_57_1_r : _tagMuxOut_T_111_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_1 = 6'h3a == index ? tagArrayWire_58_1_r : _tagMuxOut_T_113_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_1 = 6'h3b == index ? tagArrayWire_59_1_r : _tagMuxOut_T_115_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_1 = 6'h3c == index ? tagArrayWire_60_1_r : _tagMuxOut_T_117_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_1 = 6'h3d == index ? tagArrayWire_61_1_r : _tagMuxOut_T_119_1; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_1 = 6'h3e == index ? tagArrayWire_62_1_r : _tagMuxOut_T_121_1; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_1 = 6'h3f == index ? tagArrayWire_63_1_r : _tagMuxOut_T_123_1; // @[Mux.scala 80:57]
  wire  hitArray_1 = vMuxOut_1 & tagMuxOut_1 == tag; // @[Cache.scala 243:60]
  reg  vArrayWire_63_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_2_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_2_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_2 = 6'h1 == index ? vArrayWire_1_2_r : vArrayWire_0_2_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_2 = 6'h2 == index ? vArrayWire_2_2_r : _vMuxOut_T_1_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_2 = 6'h3 == index ? vArrayWire_3_2_r : _vMuxOut_T_3_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_2 = 6'h4 == index ? vArrayWire_4_2_r : _vMuxOut_T_5_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_2 = 6'h5 == index ? vArrayWire_5_2_r : _vMuxOut_T_7_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_2 = 6'h6 == index ? vArrayWire_6_2_r : _vMuxOut_T_9_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_2 = 6'h7 == index ? vArrayWire_7_2_r : _vMuxOut_T_11_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_2 = 6'h8 == index ? vArrayWire_8_2_r : _vMuxOut_T_13_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_2 = 6'h9 == index ? vArrayWire_9_2_r : _vMuxOut_T_15_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_2 = 6'ha == index ? vArrayWire_10_2_r : _vMuxOut_T_17_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_2 = 6'hb == index ? vArrayWire_11_2_r : _vMuxOut_T_19_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_2 = 6'hc == index ? vArrayWire_12_2_r : _vMuxOut_T_21_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_2 = 6'hd == index ? vArrayWire_13_2_r : _vMuxOut_T_23_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_2 = 6'he == index ? vArrayWire_14_2_r : _vMuxOut_T_25_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_2 = 6'hf == index ? vArrayWire_15_2_r : _vMuxOut_T_27_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_2 = 6'h10 == index ? vArrayWire_16_2_r : _vMuxOut_T_29_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_2 = 6'h11 == index ? vArrayWire_17_2_r : _vMuxOut_T_31_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_2 = 6'h12 == index ? vArrayWire_18_2_r : _vMuxOut_T_33_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_2 = 6'h13 == index ? vArrayWire_19_2_r : _vMuxOut_T_35_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_2 = 6'h14 == index ? vArrayWire_20_2_r : _vMuxOut_T_37_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_2 = 6'h15 == index ? vArrayWire_21_2_r : _vMuxOut_T_39_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_2 = 6'h16 == index ? vArrayWire_22_2_r : _vMuxOut_T_41_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_2 = 6'h17 == index ? vArrayWire_23_2_r : _vMuxOut_T_43_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_2 = 6'h18 == index ? vArrayWire_24_2_r : _vMuxOut_T_45_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_2 = 6'h19 == index ? vArrayWire_25_2_r : _vMuxOut_T_47_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_2 = 6'h1a == index ? vArrayWire_26_2_r : _vMuxOut_T_49_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_2 = 6'h1b == index ? vArrayWire_27_2_r : _vMuxOut_T_51_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_2 = 6'h1c == index ? vArrayWire_28_2_r : _vMuxOut_T_53_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_2 = 6'h1d == index ? vArrayWire_29_2_r : _vMuxOut_T_55_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_2 = 6'h1e == index ? vArrayWire_30_2_r : _vMuxOut_T_57_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_2 = 6'h1f == index ? vArrayWire_31_2_r : _vMuxOut_T_59_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_2 = 6'h20 == index ? vArrayWire_32_2_r : _vMuxOut_T_61_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_2 = 6'h21 == index ? vArrayWire_33_2_r : _vMuxOut_T_63_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_2 = 6'h22 == index ? vArrayWire_34_2_r : _vMuxOut_T_65_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_2 = 6'h23 == index ? vArrayWire_35_2_r : _vMuxOut_T_67_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_2 = 6'h24 == index ? vArrayWire_36_2_r : _vMuxOut_T_69_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_2 = 6'h25 == index ? vArrayWire_37_2_r : _vMuxOut_T_71_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_2 = 6'h26 == index ? vArrayWire_38_2_r : _vMuxOut_T_73_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_2 = 6'h27 == index ? vArrayWire_39_2_r : _vMuxOut_T_75_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_2 = 6'h28 == index ? vArrayWire_40_2_r : _vMuxOut_T_77_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_2 = 6'h29 == index ? vArrayWire_41_2_r : _vMuxOut_T_79_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_2 = 6'h2a == index ? vArrayWire_42_2_r : _vMuxOut_T_81_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_2 = 6'h2b == index ? vArrayWire_43_2_r : _vMuxOut_T_83_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_2 = 6'h2c == index ? vArrayWire_44_2_r : _vMuxOut_T_85_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_2 = 6'h2d == index ? vArrayWire_45_2_r : _vMuxOut_T_87_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_2 = 6'h2e == index ? vArrayWire_46_2_r : _vMuxOut_T_89_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_2 = 6'h2f == index ? vArrayWire_47_2_r : _vMuxOut_T_91_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_2 = 6'h30 == index ? vArrayWire_48_2_r : _vMuxOut_T_93_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_2 = 6'h31 == index ? vArrayWire_49_2_r : _vMuxOut_T_95_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_2 = 6'h32 == index ? vArrayWire_50_2_r : _vMuxOut_T_97_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_2 = 6'h33 == index ? vArrayWire_51_2_r : _vMuxOut_T_99_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_2 = 6'h34 == index ? vArrayWire_52_2_r : _vMuxOut_T_101_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_2 = 6'h35 == index ? vArrayWire_53_2_r : _vMuxOut_T_103_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_2 = 6'h36 == index ? vArrayWire_54_2_r : _vMuxOut_T_105_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_2 = 6'h37 == index ? vArrayWire_55_2_r : _vMuxOut_T_107_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_2 = 6'h38 == index ? vArrayWire_56_2_r : _vMuxOut_T_109_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_2 = 6'h39 == index ? vArrayWire_57_2_r : _vMuxOut_T_111_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_2 = 6'h3a == index ? vArrayWire_58_2_r : _vMuxOut_T_113_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_2 = 6'h3b == index ? vArrayWire_59_2_r : _vMuxOut_T_115_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_2 = 6'h3c == index ? vArrayWire_60_2_r : _vMuxOut_T_117_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_2 = 6'h3d == index ? vArrayWire_61_2_r : _vMuxOut_T_119_2; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_2 = 6'h3e == index ? vArrayWire_62_2_r : _vMuxOut_T_121_2; // @[Mux.scala 80:57]
  wire  vMuxOut_2 = 6'h3f == index ? vArrayWire_63_2_r : _vMuxOut_T_123_2; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_2_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_2_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_2 = 6'h1 == index ? tagArrayWire_1_2_r : tagArrayWire_0_2_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_2 = 6'h2 == index ? tagArrayWire_2_2_r : _tagMuxOut_T_1_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_2 = 6'h3 == index ? tagArrayWire_3_2_r : _tagMuxOut_T_3_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_2 = 6'h4 == index ? tagArrayWire_4_2_r : _tagMuxOut_T_5_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_2 = 6'h5 == index ? tagArrayWire_5_2_r : _tagMuxOut_T_7_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_2 = 6'h6 == index ? tagArrayWire_6_2_r : _tagMuxOut_T_9_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_2 = 6'h7 == index ? tagArrayWire_7_2_r : _tagMuxOut_T_11_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_2 = 6'h8 == index ? tagArrayWire_8_2_r : _tagMuxOut_T_13_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_2 = 6'h9 == index ? tagArrayWire_9_2_r : _tagMuxOut_T_15_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_2 = 6'ha == index ? tagArrayWire_10_2_r : _tagMuxOut_T_17_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_2 = 6'hb == index ? tagArrayWire_11_2_r : _tagMuxOut_T_19_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_2 = 6'hc == index ? tagArrayWire_12_2_r : _tagMuxOut_T_21_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_2 = 6'hd == index ? tagArrayWire_13_2_r : _tagMuxOut_T_23_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_2 = 6'he == index ? tagArrayWire_14_2_r : _tagMuxOut_T_25_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_2 = 6'hf == index ? tagArrayWire_15_2_r : _tagMuxOut_T_27_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_2 = 6'h10 == index ? tagArrayWire_16_2_r : _tagMuxOut_T_29_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_2 = 6'h11 == index ? tagArrayWire_17_2_r : _tagMuxOut_T_31_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_2 = 6'h12 == index ? tagArrayWire_18_2_r : _tagMuxOut_T_33_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_2 = 6'h13 == index ? tagArrayWire_19_2_r : _tagMuxOut_T_35_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_2 = 6'h14 == index ? tagArrayWire_20_2_r : _tagMuxOut_T_37_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_2 = 6'h15 == index ? tagArrayWire_21_2_r : _tagMuxOut_T_39_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_2 = 6'h16 == index ? tagArrayWire_22_2_r : _tagMuxOut_T_41_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_2 = 6'h17 == index ? tagArrayWire_23_2_r : _tagMuxOut_T_43_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_2 = 6'h18 == index ? tagArrayWire_24_2_r : _tagMuxOut_T_45_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_2 = 6'h19 == index ? tagArrayWire_25_2_r : _tagMuxOut_T_47_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_2 = 6'h1a == index ? tagArrayWire_26_2_r : _tagMuxOut_T_49_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_2 = 6'h1b == index ? tagArrayWire_27_2_r : _tagMuxOut_T_51_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_2 = 6'h1c == index ? tagArrayWire_28_2_r : _tagMuxOut_T_53_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_2 = 6'h1d == index ? tagArrayWire_29_2_r : _tagMuxOut_T_55_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_2 = 6'h1e == index ? tagArrayWire_30_2_r : _tagMuxOut_T_57_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_2 = 6'h1f == index ? tagArrayWire_31_2_r : _tagMuxOut_T_59_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_2 = 6'h20 == index ? tagArrayWire_32_2_r : _tagMuxOut_T_61_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_2 = 6'h21 == index ? tagArrayWire_33_2_r : _tagMuxOut_T_63_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_2 = 6'h22 == index ? tagArrayWire_34_2_r : _tagMuxOut_T_65_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_2 = 6'h23 == index ? tagArrayWire_35_2_r : _tagMuxOut_T_67_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_2 = 6'h24 == index ? tagArrayWire_36_2_r : _tagMuxOut_T_69_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_2 = 6'h25 == index ? tagArrayWire_37_2_r : _tagMuxOut_T_71_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_2 = 6'h26 == index ? tagArrayWire_38_2_r : _tagMuxOut_T_73_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_2 = 6'h27 == index ? tagArrayWire_39_2_r : _tagMuxOut_T_75_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_2 = 6'h28 == index ? tagArrayWire_40_2_r : _tagMuxOut_T_77_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_2 = 6'h29 == index ? tagArrayWire_41_2_r : _tagMuxOut_T_79_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_2 = 6'h2a == index ? tagArrayWire_42_2_r : _tagMuxOut_T_81_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_2 = 6'h2b == index ? tagArrayWire_43_2_r : _tagMuxOut_T_83_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_2 = 6'h2c == index ? tagArrayWire_44_2_r : _tagMuxOut_T_85_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_2 = 6'h2d == index ? tagArrayWire_45_2_r : _tagMuxOut_T_87_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_2 = 6'h2e == index ? tagArrayWire_46_2_r : _tagMuxOut_T_89_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_2 = 6'h2f == index ? tagArrayWire_47_2_r : _tagMuxOut_T_91_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_2 = 6'h30 == index ? tagArrayWire_48_2_r : _tagMuxOut_T_93_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_2 = 6'h31 == index ? tagArrayWire_49_2_r : _tagMuxOut_T_95_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_2 = 6'h32 == index ? tagArrayWire_50_2_r : _tagMuxOut_T_97_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_2 = 6'h33 == index ? tagArrayWire_51_2_r : _tagMuxOut_T_99_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_2 = 6'h34 == index ? tagArrayWire_52_2_r : _tagMuxOut_T_101_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_2 = 6'h35 == index ? tagArrayWire_53_2_r : _tagMuxOut_T_103_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_2 = 6'h36 == index ? tagArrayWire_54_2_r : _tagMuxOut_T_105_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_2 = 6'h37 == index ? tagArrayWire_55_2_r : _tagMuxOut_T_107_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_2 = 6'h38 == index ? tagArrayWire_56_2_r : _tagMuxOut_T_109_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_2 = 6'h39 == index ? tagArrayWire_57_2_r : _tagMuxOut_T_111_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_2 = 6'h3a == index ? tagArrayWire_58_2_r : _tagMuxOut_T_113_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_2 = 6'h3b == index ? tagArrayWire_59_2_r : _tagMuxOut_T_115_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_2 = 6'h3c == index ? tagArrayWire_60_2_r : _tagMuxOut_T_117_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_2 = 6'h3d == index ? tagArrayWire_61_2_r : _tagMuxOut_T_119_2; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_2 = 6'h3e == index ? tagArrayWire_62_2_r : _tagMuxOut_T_121_2; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_2 = 6'h3f == index ? tagArrayWire_63_2_r : _tagMuxOut_T_123_2; // @[Mux.scala 80:57]
  wire  hitArray_2 = vMuxOut_2 & tagMuxOut_2 == tag; // @[Cache.scala 243:60]
  reg  vArrayWire_63_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_62_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_61_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_60_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_59_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_58_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_57_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_56_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_55_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_54_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_53_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_52_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_51_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_50_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_49_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_48_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_47_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_46_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_45_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_44_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_43_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_42_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_41_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_40_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_39_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_38_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_37_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_36_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_35_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_34_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_33_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_32_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_31_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_30_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_29_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_28_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_27_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_26_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_25_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_24_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_23_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_22_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_21_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_20_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_19_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_18_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_17_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_16_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_15_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_14_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_13_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_12_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_11_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_10_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_9_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_8_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_7_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_6_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_5_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_4_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_3_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_2_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_1_3_r; // @[Reg.scala 27:20]
  reg  vArrayWire_0_3_r; // @[Reg.scala 27:20]
  wire  _vMuxOut_T_1_3 = 6'h1 == index ? vArrayWire_1_3_r : vArrayWire_0_3_r; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_3_3 = 6'h2 == index ? vArrayWire_2_3_r : _vMuxOut_T_1_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_5_3 = 6'h3 == index ? vArrayWire_3_3_r : _vMuxOut_T_3_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_7_3 = 6'h4 == index ? vArrayWire_4_3_r : _vMuxOut_T_5_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_9_3 = 6'h5 == index ? vArrayWire_5_3_r : _vMuxOut_T_7_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_11_3 = 6'h6 == index ? vArrayWire_6_3_r : _vMuxOut_T_9_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_13_3 = 6'h7 == index ? vArrayWire_7_3_r : _vMuxOut_T_11_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_15_3 = 6'h8 == index ? vArrayWire_8_3_r : _vMuxOut_T_13_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_17_3 = 6'h9 == index ? vArrayWire_9_3_r : _vMuxOut_T_15_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_19_3 = 6'ha == index ? vArrayWire_10_3_r : _vMuxOut_T_17_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_21_3 = 6'hb == index ? vArrayWire_11_3_r : _vMuxOut_T_19_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_23_3 = 6'hc == index ? vArrayWire_12_3_r : _vMuxOut_T_21_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_25_3 = 6'hd == index ? vArrayWire_13_3_r : _vMuxOut_T_23_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_27_3 = 6'he == index ? vArrayWire_14_3_r : _vMuxOut_T_25_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_29_3 = 6'hf == index ? vArrayWire_15_3_r : _vMuxOut_T_27_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_31_3 = 6'h10 == index ? vArrayWire_16_3_r : _vMuxOut_T_29_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_33_3 = 6'h11 == index ? vArrayWire_17_3_r : _vMuxOut_T_31_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_35_3 = 6'h12 == index ? vArrayWire_18_3_r : _vMuxOut_T_33_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_37_3 = 6'h13 == index ? vArrayWire_19_3_r : _vMuxOut_T_35_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_39_3 = 6'h14 == index ? vArrayWire_20_3_r : _vMuxOut_T_37_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_41_3 = 6'h15 == index ? vArrayWire_21_3_r : _vMuxOut_T_39_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_43_3 = 6'h16 == index ? vArrayWire_22_3_r : _vMuxOut_T_41_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_45_3 = 6'h17 == index ? vArrayWire_23_3_r : _vMuxOut_T_43_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_47_3 = 6'h18 == index ? vArrayWire_24_3_r : _vMuxOut_T_45_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_49_3 = 6'h19 == index ? vArrayWire_25_3_r : _vMuxOut_T_47_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_51_3 = 6'h1a == index ? vArrayWire_26_3_r : _vMuxOut_T_49_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_53_3 = 6'h1b == index ? vArrayWire_27_3_r : _vMuxOut_T_51_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_55_3 = 6'h1c == index ? vArrayWire_28_3_r : _vMuxOut_T_53_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_57_3 = 6'h1d == index ? vArrayWire_29_3_r : _vMuxOut_T_55_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_59_3 = 6'h1e == index ? vArrayWire_30_3_r : _vMuxOut_T_57_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_61_3 = 6'h1f == index ? vArrayWire_31_3_r : _vMuxOut_T_59_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_63_3 = 6'h20 == index ? vArrayWire_32_3_r : _vMuxOut_T_61_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_65_3 = 6'h21 == index ? vArrayWire_33_3_r : _vMuxOut_T_63_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_67_3 = 6'h22 == index ? vArrayWire_34_3_r : _vMuxOut_T_65_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_69_3 = 6'h23 == index ? vArrayWire_35_3_r : _vMuxOut_T_67_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_71_3 = 6'h24 == index ? vArrayWire_36_3_r : _vMuxOut_T_69_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_73_3 = 6'h25 == index ? vArrayWire_37_3_r : _vMuxOut_T_71_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_75_3 = 6'h26 == index ? vArrayWire_38_3_r : _vMuxOut_T_73_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_77_3 = 6'h27 == index ? vArrayWire_39_3_r : _vMuxOut_T_75_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_79_3 = 6'h28 == index ? vArrayWire_40_3_r : _vMuxOut_T_77_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_81_3 = 6'h29 == index ? vArrayWire_41_3_r : _vMuxOut_T_79_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_83_3 = 6'h2a == index ? vArrayWire_42_3_r : _vMuxOut_T_81_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_85_3 = 6'h2b == index ? vArrayWire_43_3_r : _vMuxOut_T_83_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_87_3 = 6'h2c == index ? vArrayWire_44_3_r : _vMuxOut_T_85_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_89_3 = 6'h2d == index ? vArrayWire_45_3_r : _vMuxOut_T_87_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_91_3 = 6'h2e == index ? vArrayWire_46_3_r : _vMuxOut_T_89_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_93_3 = 6'h2f == index ? vArrayWire_47_3_r : _vMuxOut_T_91_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_95_3 = 6'h30 == index ? vArrayWire_48_3_r : _vMuxOut_T_93_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_97_3 = 6'h31 == index ? vArrayWire_49_3_r : _vMuxOut_T_95_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_99_3 = 6'h32 == index ? vArrayWire_50_3_r : _vMuxOut_T_97_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_101_3 = 6'h33 == index ? vArrayWire_51_3_r : _vMuxOut_T_99_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_103_3 = 6'h34 == index ? vArrayWire_52_3_r : _vMuxOut_T_101_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_105_3 = 6'h35 == index ? vArrayWire_53_3_r : _vMuxOut_T_103_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_107_3 = 6'h36 == index ? vArrayWire_54_3_r : _vMuxOut_T_105_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_109_3 = 6'h37 == index ? vArrayWire_55_3_r : _vMuxOut_T_107_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_111_3 = 6'h38 == index ? vArrayWire_56_3_r : _vMuxOut_T_109_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_113_3 = 6'h39 == index ? vArrayWire_57_3_r : _vMuxOut_T_111_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_115_3 = 6'h3a == index ? vArrayWire_58_3_r : _vMuxOut_T_113_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_117_3 = 6'h3b == index ? vArrayWire_59_3_r : _vMuxOut_T_115_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_119_3 = 6'h3c == index ? vArrayWire_60_3_r : _vMuxOut_T_117_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_121_3 = 6'h3d == index ? vArrayWire_61_3_r : _vMuxOut_T_119_3; // @[Mux.scala 80:57]
  wire  _vMuxOut_T_123_3 = 6'h3e == index ? vArrayWire_62_3_r : _vMuxOut_T_121_3; // @[Mux.scala 80:57]
  wire  vMuxOut_3 = 6'h3f == index ? vArrayWire_63_3_r : _vMuxOut_T_123_3; // @[Mux.scala 80:57]
  reg [21:0] tagArrayWire_63_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_62_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_61_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_60_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_59_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_58_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_57_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_56_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_55_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_54_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_53_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_52_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_51_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_50_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_49_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_48_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_47_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_46_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_45_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_44_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_43_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_42_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_41_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_40_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_39_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_38_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_37_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_36_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_35_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_34_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_33_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_32_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_31_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_30_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_29_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_28_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_27_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_26_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_25_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_24_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_23_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_22_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_21_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_20_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_19_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_18_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_17_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_16_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_15_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_14_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_13_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_12_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_11_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_10_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_9_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_8_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_7_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_6_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_5_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_4_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_3_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_2_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_1_3_r; // @[Reg.scala 27:20]
  reg [21:0] tagArrayWire_0_3_r; // @[Reg.scala 27:20]
  wire [21:0] _tagMuxOut_T_1_3 = 6'h1 == index ? tagArrayWire_1_3_r : tagArrayWire_0_3_r; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_3_3 = 6'h2 == index ? tagArrayWire_2_3_r : _tagMuxOut_T_1_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_5_3 = 6'h3 == index ? tagArrayWire_3_3_r : _tagMuxOut_T_3_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_7_3 = 6'h4 == index ? tagArrayWire_4_3_r : _tagMuxOut_T_5_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_9_3 = 6'h5 == index ? tagArrayWire_5_3_r : _tagMuxOut_T_7_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_11_3 = 6'h6 == index ? tagArrayWire_6_3_r : _tagMuxOut_T_9_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_13_3 = 6'h7 == index ? tagArrayWire_7_3_r : _tagMuxOut_T_11_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_15_3 = 6'h8 == index ? tagArrayWire_8_3_r : _tagMuxOut_T_13_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_17_3 = 6'h9 == index ? tagArrayWire_9_3_r : _tagMuxOut_T_15_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_19_3 = 6'ha == index ? tagArrayWire_10_3_r : _tagMuxOut_T_17_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_21_3 = 6'hb == index ? tagArrayWire_11_3_r : _tagMuxOut_T_19_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_23_3 = 6'hc == index ? tagArrayWire_12_3_r : _tagMuxOut_T_21_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_25_3 = 6'hd == index ? tagArrayWire_13_3_r : _tagMuxOut_T_23_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_27_3 = 6'he == index ? tagArrayWire_14_3_r : _tagMuxOut_T_25_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_29_3 = 6'hf == index ? tagArrayWire_15_3_r : _tagMuxOut_T_27_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_31_3 = 6'h10 == index ? tagArrayWire_16_3_r : _tagMuxOut_T_29_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_33_3 = 6'h11 == index ? tagArrayWire_17_3_r : _tagMuxOut_T_31_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_35_3 = 6'h12 == index ? tagArrayWire_18_3_r : _tagMuxOut_T_33_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_37_3 = 6'h13 == index ? tagArrayWire_19_3_r : _tagMuxOut_T_35_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_39_3 = 6'h14 == index ? tagArrayWire_20_3_r : _tagMuxOut_T_37_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_41_3 = 6'h15 == index ? tagArrayWire_21_3_r : _tagMuxOut_T_39_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_43_3 = 6'h16 == index ? tagArrayWire_22_3_r : _tagMuxOut_T_41_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_45_3 = 6'h17 == index ? tagArrayWire_23_3_r : _tagMuxOut_T_43_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_47_3 = 6'h18 == index ? tagArrayWire_24_3_r : _tagMuxOut_T_45_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_49_3 = 6'h19 == index ? tagArrayWire_25_3_r : _tagMuxOut_T_47_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_51_3 = 6'h1a == index ? tagArrayWire_26_3_r : _tagMuxOut_T_49_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_53_3 = 6'h1b == index ? tagArrayWire_27_3_r : _tagMuxOut_T_51_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_55_3 = 6'h1c == index ? tagArrayWire_28_3_r : _tagMuxOut_T_53_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_57_3 = 6'h1d == index ? tagArrayWire_29_3_r : _tagMuxOut_T_55_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_59_3 = 6'h1e == index ? tagArrayWire_30_3_r : _tagMuxOut_T_57_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_61_3 = 6'h1f == index ? tagArrayWire_31_3_r : _tagMuxOut_T_59_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_63_3 = 6'h20 == index ? tagArrayWire_32_3_r : _tagMuxOut_T_61_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_65_3 = 6'h21 == index ? tagArrayWire_33_3_r : _tagMuxOut_T_63_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_67_3 = 6'h22 == index ? tagArrayWire_34_3_r : _tagMuxOut_T_65_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_69_3 = 6'h23 == index ? tagArrayWire_35_3_r : _tagMuxOut_T_67_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_71_3 = 6'h24 == index ? tagArrayWire_36_3_r : _tagMuxOut_T_69_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_73_3 = 6'h25 == index ? tagArrayWire_37_3_r : _tagMuxOut_T_71_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_75_3 = 6'h26 == index ? tagArrayWire_38_3_r : _tagMuxOut_T_73_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_77_3 = 6'h27 == index ? tagArrayWire_39_3_r : _tagMuxOut_T_75_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_79_3 = 6'h28 == index ? tagArrayWire_40_3_r : _tagMuxOut_T_77_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_81_3 = 6'h29 == index ? tagArrayWire_41_3_r : _tagMuxOut_T_79_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_83_3 = 6'h2a == index ? tagArrayWire_42_3_r : _tagMuxOut_T_81_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_85_3 = 6'h2b == index ? tagArrayWire_43_3_r : _tagMuxOut_T_83_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_87_3 = 6'h2c == index ? tagArrayWire_44_3_r : _tagMuxOut_T_85_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_89_3 = 6'h2d == index ? tagArrayWire_45_3_r : _tagMuxOut_T_87_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_91_3 = 6'h2e == index ? tagArrayWire_46_3_r : _tagMuxOut_T_89_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_93_3 = 6'h2f == index ? tagArrayWire_47_3_r : _tagMuxOut_T_91_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_95_3 = 6'h30 == index ? tagArrayWire_48_3_r : _tagMuxOut_T_93_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_97_3 = 6'h31 == index ? tagArrayWire_49_3_r : _tagMuxOut_T_95_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_99_3 = 6'h32 == index ? tagArrayWire_50_3_r : _tagMuxOut_T_97_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_101_3 = 6'h33 == index ? tagArrayWire_51_3_r : _tagMuxOut_T_99_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_103_3 = 6'h34 == index ? tagArrayWire_52_3_r : _tagMuxOut_T_101_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_105_3 = 6'h35 == index ? tagArrayWire_53_3_r : _tagMuxOut_T_103_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_107_3 = 6'h36 == index ? tagArrayWire_54_3_r : _tagMuxOut_T_105_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_109_3 = 6'h37 == index ? tagArrayWire_55_3_r : _tagMuxOut_T_107_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_111_3 = 6'h38 == index ? tagArrayWire_56_3_r : _tagMuxOut_T_109_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_113_3 = 6'h39 == index ? tagArrayWire_57_3_r : _tagMuxOut_T_111_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_115_3 = 6'h3a == index ? tagArrayWire_58_3_r : _tagMuxOut_T_113_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_117_3 = 6'h3b == index ? tagArrayWire_59_3_r : _tagMuxOut_T_115_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_119_3 = 6'h3c == index ? tagArrayWire_60_3_r : _tagMuxOut_T_117_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_121_3 = 6'h3d == index ? tagArrayWire_61_3_r : _tagMuxOut_T_119_3; // @[Mux.scala 80:57]
  wire [21:0] _tagMuxOut_T_123_3 = 6'h3e == index ? tagArrayWire_62_3_r : _tagMuxOut_T_121_3; // @[Mux.scala 80:57]
  wire [21:0] tagMuxOut_3 = 6'h3f == index ? tagArrayWire_63_3_r : _tagMuxOut_T_123_3; // @[Mux.scala 80:57]
  wire  hitArray_3 = vMuxOut_3 & tagMuxOut_3 == tag; // @[Cache.scala 243:60]
  wire  hit = hitArray_0 | hitArray_1 | hitArray_2 | hitArray_3; // @[Cache.scala 244:49]
  wire [1:0] _IdleMux_T_2 = hit ? 2'h0 : 2'h1; // @[Cache.scala 186:10]
  wire [1:0] _IdleMux_T_3 = io_cacheIn_wen ? 2'h2 : _IdleMux_T_2; // @[Cache.scala 183:8]
  wire [1:0] IdleMux = _IdleMux_T_1 ? _IdleMux_T_3 : 2'h0; // @[Cache.scala 181:20]
  wire [1:0] missMux = io_cacheOut_r_last_i ? 2'h0 : 2'h1; // @[Cache.scala 194:20]
  wire [1:0] _writeMux_T = io_block ? 2'h3 : 2'h0; // @[Cache.scala 197:8]
  wire  isIdle = cacheState == 2'h0; // @[Cache.scala 214:27]
  wire  isMiss = cacheState == 2'h1; // @[Cache.scala 215:27]
  wire  isWrite = cacheState == 2'h2; // @[Cache.scala 216:28]
  wire  isBlock = cacheState == 2'h3; // @[Cache.scala 217:28]
  wire [127:0] _waysel_T = hitArray_0 ? io_SRAMIO_0_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_1 = hitArray_1 ? io_SRAMIO_1_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_2 = hitArray_2 ? io_SRAMIO_2_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_3 = hitArray_3 ? io_SRAMIO_3_rdata : 128'h0; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_4 = _waysel_T | _waysel_T_1; // @[Mux.scala 27:72]
  wire [127:0] _waysel_T_5 = _waysel_T_4 | _waysel_T_2; // @[Mux.scala 27:72]
  wire [127:0] waysel = _waysel_T_5 | _waysel_T_3; // @[Mux.scala 27:72]
  reg [1:0] selArrayWire_1_r; // @[Reg.scala 27:20]
  reg [1:0] selArrayWire_0_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_1 = 6'h1 == index ? selArrayWire_1_r : selArrayWire_0_r; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_2_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_3 = 6'h2 == index ? selArrayWire_2_r : _sramSel_T_1; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_3_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_5 = 6'h3 == index ? selArrayWire_3_r : _sramSel_T_3; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_4_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_7 = 6'h4 == index ? selArrayWire_4_r : _sramSel_T_5; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_5_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_9 = 6'h5 == index ? selArrayWire_5_r : _sramSel_T_7; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_6_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_11 = 6'h6 == index ? selArrayWire_6_r : _sramSel_T_9; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_7_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_13 = 6'h7 == index ? selArrayWire_7_r : _sramSel_T_11; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_8_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_15 = 6'h8 == index ? selArrayWire_8_r : _sramSel_T_13; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_9_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_17 = 6'h9 == index ? selArrayWire_9_r : _sramSel_T_15; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_10_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_19 = 6'ha == index ? selArrayWire_10_r : _sramSel_T_17; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_11_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_21 = 6'hb == index ? selArrayWire_11_r : _sramSel_T_19; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_12_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_23 = 6'hc == index ? selArrayWire_12_r : _sramSel_T_21; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_13_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_25 = 6'hd == index ? selArrayWire_13_r : _sramSel_T_23; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_14_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_27 = 6'he == index ? selArrayWire_14_r : _sramSel_T_25; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_15_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_29 = 6'hf == index ? selArrayWire_15_r : _sramSel_T_27; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_16_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_31 = 6'h10 == index ? selArrayWire_16_r : _sramSel_T_29; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_17_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_33 = 6'h11 == index ? selArrayWire_17_r : _sramSel_T_31; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_18_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_35 = 6'h12 == index ? selArrayWire_18_r : _sramSel_T_33; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_19_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_37 = 6'h13 == index ? selArrayWire_19_r : _sramSel_T_35; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_20_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_39 = 6'h14 == index ? selArrayWire_20_r : _sramSel_T_37; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_21_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_41 = 6'h15 == index ? selArrayWire_21_r : _sramSel_T_39; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_22_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_43 = 6'h16 == index ? selArrayWire_22_r : _sramSel_T_41; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_23_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_45 = 6'h17 == index ? selArrayWire_23_r : _sramSel_T_43; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_24_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_47 = 6'h18 == index ? selArrayWire_24_r : _sramSel_T_45; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_25_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_49 = 6'h19 == index ? selArrayWire_25_r : _sramSel_T_47; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_26_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_51 = 6'h1a == index ? selArrayWire_26_r : _sramSel_T_49; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_27_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_53 = 6'h1b == index ? selArrayWire_27_r : _sramSel_T_51; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_28_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_55 = 6'h1c == index ? selArrayWire_28_r : _sramSel_T_53; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_29_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_57 = 6'h1d == index ? selArrayWire_29_r : _sramSel_T_55; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_30_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_59 = 6'h1e == index ? selArrayWire_30_r : _sramSel_T_57; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_31_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_61 = 6'h1f == index ? selArrayWire_31_r : _sramSel_T_59; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_32_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_63 = 6'h20 == index ? selArrayWire_32_r : _sramSel_T_61; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_33_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_65 = 6'h21 == index ? selArrayWire_33_r : _sramSel_T_63; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_34_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_67 = 6'h22 == index ? selArrayWire_34_r : _sramSel_T_65; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_35_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_69 = 6'h23 == index ? selArrayWire_35_r : _sramSel_T_67; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_36_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_71 = 6'h24 == index ? selArrayWire_36_r : _sramSel_T_69; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_37_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_73 = 6'h25 == index ? selArrayWire_37_r : _sramSel_T_71; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_38_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_75 = 6'h26 == index ? selArrayWire_38_r : _sramSel_T_73; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_39_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_77 = 6'h27 == index ? selArrayWire_39_r : _sramSel_T_75; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_40_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_79 = 6'h28 == index ? selArrayWire_40_r : _sramSel_T_77; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_41_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_81 = 6'h29 == index ? selArrayWire_41_r : _sramSel_T_79; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_42_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_83 = 6'h2a == index ? selArrayWire_42_r : _sramSel_T_81; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_43_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_85 = 6'h2b == index ? selArrayWire_43_r : _sramSel_T_83; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_44_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_87 = 6'h2c == index ? selArrayWire_44_r : _sramSel_T_85; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_45_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_89 = 6'h2d == index ? selArrayWire_45_r : _sramSel_T_87; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_46_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_91 = 6'h2e == index ? selArrayWire_46_r : _sramSel_T_89; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_47_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_93 = 6'h2f == index ? selArrayWire_47_r : _sramSel_T_91; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_48_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_95 = 6'h30 == index ? selArrayWire_48_r : _sramSel_T_93; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_49_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_97 = 6'h31 == index ? selArrayWire_49_r : _sramSel_T_95; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_50_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_99 = 6'h32 == index ? selArrayWire_50_r : _sramSel_T_97; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_51_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_101 = 6'h33 == index ? selArrayWire_51_r : _sramSel_T_99; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_52_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_103 = 6'h34 == index ? selArrayWire_52_r : _sramSel_T_101; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_53_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_105 = 6'h35 == index ? selArrayWire_53_r : _sramSel_T_103; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_54_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_107 = 6'h36 == index ? selArrayWire_54_r : _sramSel_T_105; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_55_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_109 = 6'h37 == index ? selArrayWire_55_r : _sramSel_T_107; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_56_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_111 = 6'h38 == index ? selArrayWire_56_r : _sramSel_T_109; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_57_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_113 = 6'h39 == index ? selArrayWire_57_r : _sramSel_T_111; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_58_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_115 = 6'h3a == index ? selArrayWire_58_r : _sramSel_T_113; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_59_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_117 = 6'h3b == index ? selArrayWire_59_r : _sramSel_T_115; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_60_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_119 = 6'h3c == index ? selArrayWire_60_r : _sramSel_T_117; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_61_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_121 = 6'h3d == index ? selArrayWire_61_r : _sramSel_T_119; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_62_r; // @[Reg.scala 27:20]
  wire [1:0] _sramSel_T_123 = 6'h3e == index ? selArrayWire_62_r : _sramSel_T_121; // @[Mux.scala 80:57]
  reg [1:0] selArrayWire_63_r; // @[Reg.scala 27:20]
  wire [1:0] sramSel = 6'h3f == index ? selArrayWire_63_r : _sramSel_T_123; // @[Mux.scala 80:57]
  wire [27:0] io_cacheOut_ar_addr_o_hi = io_cacheIn_addr[31:4]; // @[Cache.scala 275:48]
  wire [1:0] _selArrayWire_0_T_1 = selArrayWire_0_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_0_T_3 = io_cacheOut_r_last_i & 6'h0 == index; // @[Cache.scala 292:28]
  wire  _tagArrayWire_0_0_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_2 = _tagArrayWire_0_0_T_4 | vArrayWire_0_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_1_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_4 = _tagArrayWire_0_1_T_4 | vArrayWire_0_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_2_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_6 = _tagArrayWire_0_2_T_4 | vArrayWire_0_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_0_3_T_4 = _selArrayWire_0_T_3 & selArrayWire_0_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_8 = _tagArrayWire_0_3_T_4 | vArrayWire_0_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_1_T_1 = selArrayWire_1_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_1_T_3 = io_cacheOut_r_last_i & _vMuxOut_T; // @[Cache.scala 292:28]
  wire  _tagArrayWire_1_0_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_11 = _tagArrayWire_1_0_T_4 | vArrayWire_1_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_1_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_13 = _tagArrayWire_1_1_T_4 | vArrayWire_1_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_2_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_15 = _tagArrayWire_1_2_T_4 | vArrayWire_1_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_1_3_T_4 = _selArrayWire_1_T_3 & selArrayWire_1_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_17 = _tagArrayWire_1_3_T_4 | vArrayWire_1_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_2_T_1 = selArrayWire_2_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_2_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_2; // @[Cache.scala 292:28]
  wire  _tagArrayWire_2_0_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_20 = _tagArrayWire_2_0_T_4 | vArrayWire_2_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_1_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_22 = _tagArrayWire_2_1_T_4 | vArrayWire_2_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_2_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_24 = _tagArrayWire_2_2_T_4 | vArrayWire_2_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_2_3_T_4 = _selArrayWire_2_T_3 & selArrayWire_2_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_26 = _tagArrayWire_2_3_T_4 | vArrayWire_2_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_3_T_1 = selArrayWire_3_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_3_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_4; // @[Cache.scala 292:28]
  wire  _tagArrayWire_3_0_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_29 = _tagArrayWire_3_0_T_4 | vArrayWire_3_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_1_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_31 = _tagArrayWire_3_1_T_4 | vArrayWire_3_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_2_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_33 = _tagArrayWire_3_2_T_4 | vArrayWire_3_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_3_3_T_4 = _selArrayWire_3_T_3 & selArrayWire_3_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_35 = _tagArrayWire_3_3_T_4 | vArrayWire_3_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_4_T_1 = selArrayWire_4_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_4_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_6; // @[Cache.scala 292:28]
  wire  _tagArrayWire_4_0_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_38 = _tagArrayWire_4_0_T_4 | vArrayWire_4_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_1_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_40 = _tagArrayWire_4_1_T_4 | vArrayWire_4_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_2_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_42 = _tagArrayWire_4_2_T_4 | vArrayWire_4_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_4_3_T_4 = _selArrayWire_4_T_3 & selArrayWire_4_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_44 = _tagArrayWire_4_3_T_4 | vArrayWire_4_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_5_T_1 = selArrayWire_5_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_5_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_8; // @[Cache.scala 292:28]
  wire  _tagArrayWire_5_0_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_47 = _tagArrayWire_5_0_T_4 | vArrayWire_5_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_1_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_49 = _tagArrayWire_5_1_T_4 | vArrayWire_5_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_2_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_51 = _tagArrayWire_5_2_T_4 | vArrayWire_5_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_5_3_T_4 = _selArrayWire_5_T_3 & selArrayWire_5_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_53 = _tagArrayWire_5_3_T_4 | vArrayWire_5_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_6_T_1 = selArrayWire_6_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_6_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_10; // @[Cache.scala 292:28]
  wire  _tagArrayWire_6_0_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_56 = _tagArrayWire_6_0_T_4 | vArrayWire_6_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_1_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_58 = _tagArrayWire_6_1_T_4 | vArrayWire_6_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_2_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_60 = _tagArrayWire_6_2_T_4 | vArrayWire_6_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_6_3_T_4 = _selArrayWire_6_T_3 & selArrayWire_6_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_62 = _tagArrayWire_6_3_T_4 | vArrayWire_6_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_7_T_1 = selArrayWire_7_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_7_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_12; // @[Cache.scala 292:28]
  wire  _tagArrayWire_7_0_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_65 = _tagArrayWire_7_0_T_4 | vArrayWire_7_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_1_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_67 = _tagArrayWire_7_1_T_4 | vArrayWire_7_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_2_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_69 = _tagArrayWire_7_2_T_4 | vArrayWire_7_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_7_3_T_4 = _selArrayWire_7_T_3 & selArrayWire_7_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_71 = _tagArrayWire_7_3_T_4 | vArrayWire_7_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_8_T_1 = selArrayWire_8_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_8_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_14; // @[Cache.scala 292:28]
  wire  _tagArrayWire_8_0_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_74 = _tagArrayWire_8_0_T_4 | vArrayWire_8_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_1_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_76 = _tagArrayWire_8_1_T_4 | vArrayWire_8_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_2_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_78 = _tagArrayWire_8_2_T_4 | vArrayWire_8_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_8_3_T_4 = _selArrayWire_8_T_3 & selArrayWire_8_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_80 = _tagArrayWire_8_3_T_4 | vArrayWire_8_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_9_T_1 = selArrayWire_9_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_9_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_16; // @[Cache.scala 292:28]
  wire  _tagArrayWire_9_0_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_83 = _tagArrayWire_9_0_T_4 | vArrayWire_9_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_1_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_85 = _tagArrayWire_9_1_T_4 | vArrayWire_9_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_2_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_87 = _tagArrayWire_9_2_T_4 | vArrayWire_9_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_9_3_T_4 = _selArrayWire_9_T_3 & selArrayWire_9_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_89 = _tagArrayWire_9_3_T_4 | vArrayWire_9_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_10_T_1 = selArrayWire_10_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_10_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_18; // @[Cache.scala 292:28]
  wire  _tagArrayWire_10_0_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_92 = _tagArrayWire_10_0_T_4 | vArrayWire_10_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_1_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_94 = _tagArrayWire_10_1_T_4 | vArrayWire_10_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_2_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_96 = _tagArrayWire_10_2_T_4 | vArrayWire_10_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_10_3_T_4 = _selArrayWire_10_T_3 & selArrayWire_10_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_98 = _tagArrayWire_10_3_T_4 | vArrayWire_10_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_11_T_1 = selArrayWire_11_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_11_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_20; // @[Cache.scala 292:28]
  wire  _tagArrayWire_11_0_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_101 = _tagArrayWire_11_0_T_4 | vArrayWire_11_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_1_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_103 = _tagArrayWire_11_1_T_4 | vArrayWire_11_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_2_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_105 = _tagArrayWire_11_2_T_4 | vArrayWire_11_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_11_3_T_4 = _selArrayWire_11_T_3 & selArrayWire_11_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_107 = _tagArrayWire_11_3_T_4 | vArrayWire_11_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_12_T_1 = selArrayWire_12_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_12_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_22; // @[Cache.scala 292:28]
  wire  _tagArrayWire_12_0_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_110 = _tagArrayWire_12_0_T_4 | vArrayWire_12_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_1_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_112 = _tagArrayWire_12_1_T_4 | vArrayWire_12_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_2_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_114 = _tagArrayWire_12_2_T_4 | vArrayWire_12_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_12_3_T_4 = _selArrayWire_12_T_3 & selArrayWire_12_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_116 = _tagArrayWire_12_3_T_4 | vArrayWire_12_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_13_T_1 = selArrayWire_13_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_13_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_24; // @[Cache.scala 292:28]
  wire  _tagArrayWire_13_0_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_119 = _tagArrayWire_13_0_T_4 | vArrayWire_13_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_1_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_121 = _tagArrayWire_13_1_T_4 | vArrayWire_13_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_2_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_123 = _tagArrayWire_13_2_T_4 | vArrayWire_13_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_13_3_T_4 = _selArrayWire_13_T_3 & selArrayWire_13_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_125 = _tagArrayWire_13_3_T_4 | vArrayWire_13_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_14_T_1 = selArrayWire_14_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_14_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_26; // @[Cache.scala 292:28]
  wire  _tagArrayWire_14_0_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_128 = _tagArrayWire_14_0_T_4 | vArrayWire_14_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_1_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_130 = _tagArrayWire_14_1_T_4 | vArrayWire_14_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_2_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_132 = _tagArrayWire_14_2_T_4 | vArrayWire_14_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_14_3_T_4 = _selArrayWire_14_T_3 & selArrayWire_14_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_134 = _tagArrayWire_14_3_T_4 | vArrayWire_14_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_15_T_1 = selArrayWire_15_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_15_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_28; // @[Cache.scala 292:28]
  wire  _tagArrayWire_15_0_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_137 = _tagArrayWire_15_0_T_4 | vArrayWire_15_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_1_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_139 = _tagArrayWire_15_1_T_4 | vArrayWire_15_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_2_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_141 = _tagArrayWire_15_2_T_4 | vArrayWire_15_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_15_3_T_4 = _selArrayWire_15_T_3 & selArrayWire_15_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_143 = _tagArrayWire_15_3_T_4 | vArrayWire_15_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_16_T_1 = selArrayWire_16_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_16_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_30; // @[Cache.scala 292:28]
  wire  _tagArrayWire_16_0_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_146 = _tagArrayWire_16_0_T_4 | vArrayWire_16_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_1_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_148 = _tagArrayWire_16_1_T_4 | vArrayWire_16_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_2_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_150 = _tagArrayWire_16_2_T_4 | vArrayWire_16_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_16_3_T_4 = _selArrayWire_16_T_3 & selArrayWire_16_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_152 = _tagArrayWire_16_3_T_4 | vArrayWire_16_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_17_T_1 = selArrayWire_17_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_17_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_32; // @[Cache.scala 292:28]
  wire  _tagArrayWire_17_0_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_155 = _tagArrayWire_17_0_T_4 | vArrayWire_17_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_1_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_157 = _tagArrayWire_17_1_T_4 | vArrayWire_17_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_2_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_159 = _tagArrayWire_17_2_T_4 | vArrayWire_17_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_17_3_T_4 = _selArrayWire_17_T_3 & selArrayWire_17_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_161 = _tagArrayWire_17_3_T_4 | vArrayWire_17_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_18_T_1 = selArrayWire_18_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_18_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_34; // @[Cache.scala 292:28]
  wire  _tagArrayWire_18_0_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_164 = _tagArrayWire_18_0_T_4 | vArrayWire_18_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_1_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_166 = _tagArrayWire_18_1_T_4 | vArrayWire_18_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_2_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_168 = _tagArrayWire_18_2_T_4 | vArrayWire_18_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_18_3_T_4 = _selArrayWire_18_T_3 & selArrayWire_18_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_170 = _tagArrayWire_18_3_T_4 | vArrayWire_18_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_19_T_1 = selArrayWire_19_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_19_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_36; // @[Cache.scala 292:28]
  wire  _tagArrayWire_19_0_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_173 = _tagArrayWire_19_0_T_4 | vArrayWire_19_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_1_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_175 = _tagArrayWire_19_1_T_4 | vArrayWire_19_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_2_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_177 = _tagArrayWire_19_2_T_4 | vArrayWire_19_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_19_3_T_4 = _selArrayWire_19_T_3 & selArrayWire_19_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_179 = _tagArrayWire_19_3_T_4 | vArrayWire_19_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_20_T_1 = selArrayWire_20_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_20_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_38; // @[Cache.scala 292:28]
  wire  _tagArrayWire_20_0_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_182 = _tagArrayWire_20_0_T_4 | vArrayWire_20_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_1_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_184 = _tagArrayWire_20_1_T_4 | vArrayWire_20_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_2_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_186 = _tagArrayWire_20_2_T_4 | vArrayWire_20_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_20_3_T_4 = _selArrayWire_20_T_3 & selArrayWire_20_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_188 = _tagArrayWire_20_3_T_4 | vArrayWire_20_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_21_T_1 = selArrayWire_21_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_21_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_40; // @[Cache.scala 292:28]
  wire  _tagArrayWire_21_0_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_191 = _tagArrayWire_21_0_T_4 | vArrayWire_21_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_1_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_193 = _tagArrayWire_21_1_T_4 | vArrayWire_21_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_2_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_195 = _tagArrayWire_21_2_T_4 | vArrayWire_21_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_21_3_T_4 = _selArrayWire_21_T_3 & selArrayWire_21_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_197 = _tagArrayWire_21_3_T_4 | vArrayWire_21_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_22_T_1 = selArrayWire_22_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_22_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_42; // @[Cache.scala 292:28]
  wire  _tagArrayWire_22_0_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_200 = _tagArrayWire_22_0_T_4 | vArrayWire_22_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_1_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_202 = _tagArrayWire_22_1_T_4 | vArrayWire_22_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_2_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_204 = _tagArrayWire_22_2_T_4 | vArrayWire_22_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_22_3_T_4 = _selArrayWire_22_T_3 & selArrayWire_22_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_206 = _tagArrayWire_22_3_T_4 | vArrayWire_22_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_23_T_1 = selArrayWire_23_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_23_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_44; // @[Cache.scala 292:28]
  wire  _tagArrayWire_23_0_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_209 = _tagArrayWire_23_0_T_4 | vArrayWire_23_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_1_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_211 = _tagArrayWire_23_1_T_4 | vArrayWire_23_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_2_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_213 = _tagArrayWire_23_2_T_4 | vArrayWire_23_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_23_3_T_4 = _selArrayWire_23_T_3 & selArrayWire_23_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_215 = _tagArrayWire_23_3_T_4 | vArrayWire_23_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_24_T_1 = selArrayWire_24_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_24_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_46; // @[Cache.scala 292:28]
  wire  _tagArrayWire_24_0_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_218 = _tagArrayWire_24_0_T_4 | vArrayWire_24_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_1_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_220 = _tagArrayWire_24_1_T_4 | vArrayWire_24_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_2_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_222 = _tagArrayWire_24_2_T_4 | vArrayWire_24_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_24_3_T_4 = _selArrayWire_24_T_3 & selArrayWire_24_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_224 = _tagArrayWire_24_3_T_4 | vArrayWire_24_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_25_T_1 = selArrayWire_25_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_25_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_48; // @[Cache.scala 292:28]
  wire  _tagArrayWire_25_0_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_227 = _tagArrayWire_25_0_T_4 | vArrayWire_25_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_1_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_229 = _tagArrayWire_25_1_T_4 | vArrayWire_25_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_2_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_231 = _tagArrayWire_25_2_T_4 | vArrayWire_25_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_25_3_T_4 = _selArrayWire_25_T_3 & selArrayWire_25_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_233 = _tagArrayWire_25_3_T_4 | vArrayWire_25_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_26_T_1 = selArrayWire_26_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_26_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_50; // @[Cache.scala 292:28]
  wire  _tagArrayWire_26_0_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_236 = _tagArrayWire_26_0_T_4 | vArrayWire_26_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_1_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_238 = _tagArrayWire_26_1_T_4 | vArrayWire_26_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_2_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_240 = _tagArrayWire_26_2_T_4 | vArrayWire_26_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_26_3_T_4 = _selArrayWire_26_T_3 & selArrayWire_26_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_242 = _tagArrayWire_26_3_T_4 | vArrayWire_26_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_27_T_1 = selArrayWire_27_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_27_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_52; // @[Cache.scala 292:28]
  wire  _tagArrayWire_27_0_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_245 = _tagArrayWire_27_0_T_4 | vArrayWire_27_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_1_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_247 = _tagArrayWire_27_1_T_4 | vArrayWire_27_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_2_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_249 = _tagArrayWire_27_2_T_4 | vArrayWire_27_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_27_3_T_4 = _selArrayWire_27_T_3 & selArrayWire_27_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_251 = _tagArrayWire_27_3_T_4 | vArrayWire_27_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_28_T_1 = selArrayWire_28_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_28_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_54; // @[Cache.scala 292:28]
  wire  _tagArrayWire_28_0_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_254 = _tagArrayWire_28_0_T_4 | vArrayWire_28_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_1_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_256 = _tagArrayWire_28_1_T_4 | vArrayWire_28_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_2_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_258 = _tagArrayWire_28_2_T_4 | vArrayWire_28_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_28_3_T_4 = _selArrayWire_28_T_3 & selArrayWire_28_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_260 = _tagArrayWire_28_3_T_4 | vArrayWire_28_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_29_T_1 = selArrayWire_29_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_29_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_56; // @[Cache.scala 292:28]
  wire  _tagArrayWire_29_0_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_263 = _tagArrayWire_29_0_T_4 | vArrayWire_29_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_1_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_265 = _tagArrayWire_29_1_T_4 | vArrayWire_29_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_2_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_267 = _tagArrayWire_29_2_T_4 | vArrayWire_29_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_29_3_T_4 = _selArrayWire_29_T_3 & selArrayWire_29_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_269 = _tagArrayWire_29_3_T_4 | vArrayWire_29_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_30_T_1 = selArrayWire_30_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_30_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_58; // @[Cache.scala 292:28]
  wire  _tagArrayWire_30_0_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_272 = _tagArrayWire_30_0_T_4 | vArrayWire_30_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_1_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_274 = _tagArrayWire_30_1_T_4 | vArrayWire_30_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_2_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_276 = _tagArrayWire_30_2_T_4 | vArrayWire_30_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_30_3_T_4 = _selArrayWire_30_T_3 & selArrayWire_30_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_278 = _tagArrayWire_30_3_T_4 | vArrayWire_30_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_31_T_1 = selArrayWire_31_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_31_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_60; // @[Cache.scala 292:28]
  wire  _tagArrayWire_31_0_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_281 = _tagArrayWire_31_0_T_4 | vArrayWire_31_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_1_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_283 = _tagArrayWire_31_1_T_4 | vArrayWire_31_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_2_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_285 = _tagArrayWire_31_2_T_4 | vArrayWire_31_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_31_3_T_4 = _selArrayWire_31_T_3 & selArrayWire_31_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_287 = _tagArrayWire_31_3_T_4 | vArrayWire_31_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_32_T_1 = selArrayWire_32_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_32_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_62; // @[Cache.scala 292:28]
  wire  _tagArrayWire_32_0_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_290 = _tagArrayWire_32_0_T_4 | vArrayWire_32_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_1_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_292 = _tagArrayWire_32_1_T_4 | vArrayWire_32_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_2_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_294 = _tagArrayWire_32_2_T_4 | vArrayWire_32_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_32_3_T_4 = _selArrayWire_32_T_3 & selArrayWire_32_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_296 = _tagArrayWire_32_3_T_4 | vArrayWire_32_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_33_T_1 = selArrayWire_33_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_33_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_64; // @[Cache.scala 292:28]
  wire  _tagArrayWire_33_0_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_299 = _tagArrayWire_33_0_T_4 | vArrayWire_33_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_1_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_301 = _tagArrayWire_33_1_T_4 | vArrayWire_33_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_2_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_303 = _tagArrayWire_33_2_T_4 | vArrayWire_33_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_33_3_T_4 = _selArrayWire_33_T_3 & selArrayWire_33_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_305 = _tagArrayWire_33_3_T_4 | vArrayWire_33_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_34_T_1 = selArrayWire_34_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_34_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_66; // @[Cache.scala 292:28]
  wire  _tagArrayWire_34_0_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_308 = _tagArrayWire_34_0_T_4 | vArrayWire_34_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_1_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_310 = _tagArrayWire_34_1_T_4 | vArrayWire_34_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_2_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_312 = _tagArrayWire_34_2_T_4 | vArrayWire_34_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_34_3_T_4 = _selArrayWire_34_T_3 & selArrayWire_34_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_314 = _tagArrayWire_34_3_T_4 | vArrayWire_34_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_35_T_1 = selArrayWire_35_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_35_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_68; // @[Cache.scala 292:28]
  wire  _tagArrayWire_35_0_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_317 = _tagArrayWire_35_0_T_4 | vArrayWire_35_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_1_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_319 = _tagArrayWire_35_1_T_4 | vArrayWire_35_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_2_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_321 = _tagArrayWire_35_2_T_4 | vArrayWire_35_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_35_3_T_4 = _selArrayWire_35_T_3 & selArrayWire_35_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_323 = _tagArrayWire_35_3_T_4 | vArrayWire_35_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_36_T_1 = selArrayWire_36_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_36_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_70; // @[Cache.scala 292:28]
  wire  _tagArrayWire_36_0_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_326 = _tagArrayWire_36_0_T_4 | vArrayWire_36_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_1_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_328 = _tagArrayWire_36_1_T_4 | vArrayWire_36_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_2_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_330 = _tagArrayWire_36_2_T_4 | vArrayWire_36_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_36_3_T_4 = _selArrayWire_36_T_3 & selArrayWire_36_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_332 = _tagArrayWire_36_3_T_4 | vArrayWire_36_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_37_T_1 = selArrayWire_37_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_37_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_72; // @[Cache.scala 292:28]
  wire  _tagArrayWire_37_0_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_335 = _tagArrayWire_37_0_T_4 | vArrayWire_37_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_1_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_337 = _tagArrayWire_37_1_T_4 | vArrayWire_37_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_2_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_339 = _tagArrayWire_37_2_T_4 | vArrayWire_37_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_37_3_T_4 = _selArrayWire_37_T_3 & selArrayWire_37_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_341 = _tagArrayWire_37_3_T_4 | vArrayWire_37_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_38_T_1 = selArrayWire_38_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_38_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_74; // @[Cache.scala 292:28]
  wire  _tagArrayWire_38_0_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_344 = _tagArrayWire_38_0_T_4 | vArrayWire_38_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_1_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_346 = _tagArrayWire_38_1_T_4 | vArrayWire_38_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_2_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_348 = _tagArrayWire_38_2_T_4 | vArrayWire_38_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_38_3_T_4 = _selArrayWire_38_T_3 & selArrayWire_38_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_350 = _tagArrayWire_38_3_T_4 | vArrayWire_38_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_39_T_1 = selArrayWire_39_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_39_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_76; // @[Cache.scala 292:28]
  wire  _tagArrayWire_39_0_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_353 = _tagArrayWire_39_0_T_4 | vArrayWire_39_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_1_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_355 = _tagArrayWire_39_1_T_4 | vArrayWire_39_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_2_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_357 = _tagArrayWire_39_2_T_4 | vArrayWire_39_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_39_3_T_4 = _selArrayWire_39_T_3 & selArrayWire_39_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_359 = _tagArrayWire_39_3_T_4 | vArrayWire_39_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_40_T_1 = selArrayWire_40_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_40_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_78; // @[Cache.scala 292:28]
  wire  _tagArrayWire_40_0_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_362 = _tagArrayWire_40_0_T_4 | vArrayWire_40_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_1_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_364 = _tagArrayWire_40_1_T_4 | vArrayWire_40_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_2_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_366 = _tagArrayWire_40_2_T_4 | vArrayWire_40_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_40_3_T_4 = _selArrayWire_40_T_3 & selArrayWire_40_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_368 = _tagArrayWire_40_3_T_4 | vArrayWire_40_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_41_T_1 = selArrayWire_41_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_41_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_80; // @[Cache.scala 292:28]
  wire  _tagArrayWire_41_0_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_371 = _tagArrayWire_41_0_T_4 | vArrayWire_41_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_1_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_373 = _tagArrayWire_41_1_T_4 | vArrayWire_41_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_2_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_375 = _tagArrayWire_41_2_T_4 | vArrayWire_41_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_41_3_T_4 = _selArrayWire_41_T_3 & selArrayWire_41_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_377 = _tagArrayWire_41_3_T_4 | vArrayWire_41_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_42_T_1 = selArrayWire_42_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_42_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_82; // @[Cache.scala 292:28]
  wire  _tagArrayWire_42_0_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_380 = _tagArrayWire_42_0_T_4 | vArrayWire_42_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_1_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_382 = _tagArrayWire_42_1_T_4 | vArrayWire_42_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_2_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_384 = _tagArrayWire_42_2_T_4 | vArrayWire_42_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_42_3_T_4 = _selArrayWire_42_T_3 & selArrayWire_42_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_386 = _tagArrayWire_42_3_T_4 | vArrayWire_42_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_43_T_1 = selArrayWire_43_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_43_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_84; // @[Cache.scala 292:28]
  wire  _tagArrayWire_43_0_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_389 = _tagArrayWire_43_0_T_4 | vArrayWire_43_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_1_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_391 = _tagArrayWire_43_1_T_4 | vArrayWire_43_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_2_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_393 = _tagArrayWire_43_2_T_4 | vArrayWire_43_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_43_3_T_4 = _selArrayWire_43_T_3 & selArrayWire_43_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_395 = _tagArrayWire_43_3_T_4 | vArrayWire_43_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_44_T_1 = selArrayWire_44_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_44_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_86; // @[Cache.scala 292:28]
  wire  _tagArrayWire_44_0_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_398 = _tagArrayWire_44_0_T_4 | vArrayWire_44_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_1_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_400 = _tagArrayWire_44_1_T_4 | vArrayWire_44_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_2_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_402 = _tagArrayWire_44_2_T_4 | vArrayWire_44_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_44_3_T_4 = _selArrayWire_44_T_3 & selArrayWire_44_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_404 = _tagArrayWire_44_3_T_4 | vArrayWire_44_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_45_T_1 = selArrayWire_45_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_45_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_88; // @[Cache.scala 292:28]
  wire  _tagArrayWire_45_0_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_407 = _tagArrayWire_45_0_T_4 | vArrayWire_45_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_1_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_409 = _tagArrayWire_45_1_T_4 | vArrayWire_45_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_2_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_411 = _tagArrayWire_45_2_T_4 | vArrayWire_45_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_45_3_T_4 = _selArrayWire_45_T_3 & selArrayWire_45_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_413 = _tagArrayWire_45_3_T_4 | vArrayWire_45_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_46_T_1 = selArrayWire_46_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_46_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_90; // @[Cache.scala 292:28]
  wire  _tagArrayWire_46_0_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_416 = _tagArrayWire_46_0_T_4 | vArrayWire_46_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_1_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_418 = _tagArrayWire_46_1_T_4 | vArrayWire_46_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_2_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_420 = _tagArrayWire_46_2_T_4 | vArrayWire_46_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_46_3_T_4 = _selArrayWire_46_T_3 & selArrayWire_46_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_422 = _tagArrayWire_46_3_T_4 | vArrayWire_46_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_47_T_1 = selArrayWire_47_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_47_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_92; // @[Cache.scala 292:28]
  wire  _tagArrayWire_47_0_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_425 = _tagArrayWire_47_0_T_4 | vArrayWire_47_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_1_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_427 = _tagArrayWire_47_1_T_4 | vArrayWire_47_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_2_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_429 = _tagArrayWire_47_2_T_4 | vArrayWire_47_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_47_3_T_4 = _selArrayWire_47_T_3 & selArrayWire_47_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_431 = _tagArrayWire_47_3_T_4 | vArrayWire_47_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_48_T_1 = selArrayWire_48_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_48_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_94; // @[Cache.scala 292:28]
  wire  _tagArrayWire_48_0_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_434 = _tagArrayWire_48_0_T_4 | vArrayWire_48_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_1_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_436 = _tagArrayWire_48_1_T_4 | vArrayWire_48_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_2_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_438 = _tagArrayWire_48_2_T_4 | vArrayWire_48_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_48_3_T_4 = _selArrayWire_48_T_3 & selArrayWire_48_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_440 = _tagArrayWire_48_3_T_4 | vArrayWire_48_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_49_T_1 = selArrayWire_49_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_49_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_96; // @[Cache.scala 292:28]
  wire  _tagArrayWire_49_0_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_443 = _tagArrayWire_49_0_T_4 | vArrayWire_49_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_1_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_445 = _tagArrayWire_49_1_T_4 | vArrayWire_49_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_2_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_447 = _tagArrayWire_49_2_T_4 | vArrayWire_49_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_49_3_T_4 = _selArrayWire_49_T_3 & selArrayWire_49_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_449 = _tagArrayWire_49_3_T_4 | vArrayWire_49_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_50_T_1 = selArrayWire_50_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_50_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_98; // @[Cache.scala 292:28]
  wire  _tagArrayWire_50_0_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_452 = _tagArrayWire_50_0_T_4 | vArrayWire_50_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_1_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_454 = _tagArrayWire_50_1_T_4 | vArrayWire_50_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_2_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_456 = _tagArrayWire_50_2_T_4 | vArrayWire_50_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_50_3_T_4 = _selArrayWire_50_T_3 & selArrayWire_50_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_458 = _tagArrayWire_50_3_T_4 | vArrayWire_50_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_51_T_1 = selArrayWire_51_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_51_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_100; // @[Cache.scala 292:28]
  wire  _tagArrayWire_51_0_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_461 = _tagArrayWire_51_0_T_4 | vArrayWire_51_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_1_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_463 = _tagArrayWire_51_1_T_4 | vArrayWire_51_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_2_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_465 = _tagArrayWire_51_2_T_4 | vArrayWire_51_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_51_3_T_4 = _selArrayWire_51_T_3 & selArrayWire_51_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_467 = _tagArrayWire_51_3_T_4 | vArrayWire_51_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_52_T_1 = selArrayWire_52_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_52_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_102; // @[Cache.scala 292:28]
  wire  _tagArrayWire_52_0_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_470 = _tagArrayWire_52_0_T_4 | vArrayWire_52_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_1_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_472 = _tagArrayWire_52_1_T_4 | vArrayWire_52_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_2_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_474 = _tagArrayWire_52_2_T_4 | vArrayWire_52_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_52_3_T_4 = _selArrayWire_52_T_3 & selArrayWire_52_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_476 = _tagArrayWire_52_3_T_4 | vArrayWire_52_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_53_T_1 = selArrayWire_53_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_53_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_104; // @[Cache.scala 292:28]
  wire  _tagArrayWire_53_0_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_479 = _tagArrayWire_53_0_T_4 | vArrayWire_53_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_1_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_481 = _tagArrayWire_53_1_T_4 | vArrayWire_53_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_2_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_483 = _tagArrayWire_53_2_T_4 | vArrayWire_53_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_53_3_T_4 = _selArrayWire_53_T_3 & selArrayWire_53_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_485 = _tagArrayWire_53_3_T_4 | vArrayWire_53_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_54_T_1 = selArrayWire_54_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_54_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_106; // @[Cache.scala 292:28]
  wire  _tagArrayWire_54_0_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_488 = _tagArrayWire_54_0_T_4 | vArrayWire_54_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_1_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_490 = _tagArrayWire_54_1_T_4 | vArrayWire_54_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_2_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_492 = _tagArrayWire_54_2_T_4 | vArrayWire_54_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_54_3_T_4 = _selArrayWire_54_T_3 & selArrayWire_54_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_494 = _tagArrayWire_54_3_T_4 | vArrayWire_54_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_55_T_1 = selArrayWire_55_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_55_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_108; // @[Cache.scala 292:28]
  wire  _tagArrayWire_55_0_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_497 = _tagArrayWire_55_0_T_4 | vArrayWire_55_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_1_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_499 = _tagArrayWire_55_1_T_4 | vArrayWire_55_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_2_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_501 = _tagArrayWire_55_2_T_4 | vArrayWire_55_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_55_3_T_4 = _selArrayWire_55_T_3 & selArrayWire_55_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_503 = _tagArrayWire_55_3_T_4 | vArrayWire_55_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_56_T_1 = selArrayWire_56_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_56_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_110; // @[Cache.scala 292:28]
  wire  _tagArrayWire_56_0_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_506 = _tagArrayWire_56_0_T_4 | vArrayWire_56_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_1_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_508 = _tagArrayWire_56_1_T_4 | vArrayWire_56_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_2_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_510 = _tagArrayWire_56_2_T_4 | vArrayWire_56_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_56_3_T_4 = _selArrayWire_56_T_3 & selArrayWire_56_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_512 = _tagArrayWire_56_3_T_4 | vArrayWire_56_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_57_T_1 = selArrayWire_57_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_57_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_112; // @[Cache.scala 292:28]
  wire  _tagArrayWire_57_0_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_515 = _tagArrayWire_57_0_T_4 | vArrayWire_57_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_1_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_517 = _tagArrayWire_57_1_T_4 | vArrayWire_57_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_2_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_519 = _tagArrayWire_57_2_T_4 | vArrayWire_57_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_57_3_T_4 = _selArrayWire_57_T_3 & selArrayWire_57_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_521 = _tagArrayWire_57_3_T_4 | vArrayWire_57_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_58_T_1 = selArrayWire_58_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_58_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_114; // @[Cache.scala 292:28]
  wire  _tagArrayWire_58_0_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_524 = _tagArrayWire_58_0_T_4 | vArrayWire_58_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_1_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_526 = _tagArrayWire_58_1_T_4 | vArrayWire_58_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_2_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_528 = _tagArrayWire_58_2_T_4 | vArrayWire_58_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_58_3_T_4 = _selArrayWire_58_T_3 & selArrayWire_58_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_530 = _tagArrayWire_58_3_T_4 | vArrayWire_58_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_59_T_1 = selArrayWire_59_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_59_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_116; // @[Cache.scala 292:28]
  wire  _tagArrayWire_59_0_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_533 = _tagArrayWire_59_0_T_4 | vArrayWire_59_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_1_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_535 = _tagArrayWire_59_1_T_4 | vArrayWire_59_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_2_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_537 = _tagArrayWire_59_2_T_4 | vArrayWire_59_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_59_3_T_4 = _selArrayWire_59_T_3 & selArrayWire_59_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_539 = _tagArrayWire_59_3_T_4 | vArrayWire_59_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_60_T_1 = selArrayWire_60_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_60_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_118; // @[Cache.scala 292:28]
  wire  _tagArrayWire_60_0_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_542 = _tagArrayWire_60_0_T_4 | vArrayWire_60_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_1_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_544 = _tagArrayWire_60_1_T_4 | vArrayWire_60_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_2_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_546 = _tagArrayWire_60_2_T_4 | vArrayWire_60_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_60_3_T_4 = _selArrayWire_60_T_3 & selArrayWire_60_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_548 = _tagArrayWire_60_3_T_4 | vArrayWire_60_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_61_T_1 = selArrayWire_61_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_61_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_120; // @[Cache.scala 292:28]
  wire  _tagArrayWire_61_0_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_551 = _tagArrayWire_61_0_T_4 | vArrayWire_61_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_1_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_553 = _tagArrayWire_61_1_T_4 | vArrayWire_61_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_2_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_555 = _tagArrayWire_61_2_T_4 | vArrayWire_61_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_61_3_T_4 = _selArrayWire_61_T_3 & selArrayWire_61_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_557 = _tagArrayWire_61_3_T_4 | vArrayWire_61_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_62_T_1 = selArrayWire_62_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_62_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_122; // @[Cache.scala 292:28]
  wire  _tagArrayWire_62_0_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_560 = _tagArrayWire_62_0_T_4 | vArrayWire_62_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_1_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_562 = _tagArrayWire_62_1_T_4 | vArrayWire_62_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_2_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_564 = _tagArrayWire_62_2_T_4 | vArrayWire_62_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_62_3_T_4 = _selArrayWire_62_T_3 & selArrayWire_62_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_566 = _tagArrayWire_62_3_T_4 | vArrayWire_62_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [1:0] _selArrayWire_63_T_1 = selArrayWire_63_r + 2'h1; // @[Cache.scala 290:23]
  wire  _selArrayWire_63_T_3 = io_cacheOut_r_last_i & _vMuxOut_T_124; // @[Cache.scala 292:28]
  wire  _tagArrayWire_63_0_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h0 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_569 = _tagArrayWire_63_0_T_4 | vArrayWire_63_0_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_1_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h1 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_571 = _tagArrayWire_63_1_T_4 | vArrayWire_63_1_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_2_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h2 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_573 = _tagArrayWire_63_2_T_4 | vArrayWire_63_2_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _tagArrayWire_63_3_T_4 = _selArrayWire_63_T_3 & selArrayWire_63_r == 2'h3 & isMiss; // @[Cache.scala 295:112]
  wire  _GEN_575 = _tagArrayWire_63_3_T_4 | vArrayWire_63_3_r; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [7:0] maskWrite_0 = io_cacheIn_mask[0] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_1 = io_cacheIn_mask[1] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_2 = io_cacheIn_mask[2] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_3 = io_cacheIn_mask[3] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_4 = io_cacheIn_mask[4] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_5 = io_cacheIn_mask[5] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_6 = io_cacheIn_mask[6] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [7:0] maskWrite_7 = io_cacheIn_mask[7] ? 8'h0 : 8'hff; // @[Cache.scala 306:24]
  wire [127:0] _ramMaskWrite_T_2 = {maskWrite_7,maskWrite_6,maskWrite_5,maskWrite_4,maskWrite_3,maskWrite_2,maskWrite_1,
    maskWrite_0,64'hffffffffffffffff}; // @[Cat.scala 30:58]
  wire [127:0] _ramMaskWrite_T_4 = {64'hffffffffffffffff,maskWrite_7,maskWrite_6,maskWrite_5,maskWrite_4,maskWrite_3,
    maskWrite_2,maskWrite_1,maskWrite_0}; // @[Cat.scala 30:58]
  wire [127:0] ramMaskWrite = offset[3] ? _ramMaskWrite_T_2 : _ramMaskWrite_T_4; // @[Cache.scala 313:25]
  wire  _io_SRAMIO_0_cen_T_4 = isMiss & io_cacheOut_r_valid_i & 2'h0 == sramSel; // @[Cache.scala 341:102]
  wire [127:0] _io_SRAMIO_0_wdata_T = {io_cacheOut_r_data_i,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _io_SRAMIO_0_wdata_T_1 = {64'h0,io_cacheOut_r_data_i}; // @[Cat.scala 30:58]
  wire [127:0] _io_SRAMIO_0_wdata_T_2 = io_cacheOut_r_last_i ? _io_SRAMIO_0_wdata_T : _io_SRAMIO_0_wdata_T_1; // @[Cache.scala 346:10]
  wire [127:0] _io_SRAMIO_0_wdata_T_4 = {io_cacheIn_data_write,64'h0}; // @[Cat.scala 30:58]
  wire [127:0] _io_SRAMIO_0_wdata_T_5 = {64'h0,io_cacheIn_data_write}; // @[Cat.scala 30:58]
  wire [127:0] _io_SRAMIO_0_wdata_T_6 = offset[3] ? _io_SRAMIO_0_wdata_T_4 : _io_SRAMIO_0_wdata_T_5; // @[Cache.scala 347:10]
  wire [127:0] _io_SRAMIO_0_wmask_T_2 = io_cacheOut_r_last_i ? 128'hffffffffffffffff : 128'hffffffffffffffff0000000000000000
    ; // @[Cache.scala 351:10]
  wire  _io_SRAMIO_1_cen_T_4 = isMiss & io_cacheOut_r_valid_i & 2'h1 == sramSel; // @[Cache.scala 341:102]
  wire  _io_SRAMIO_2_cen_T_4 = isMiss & io_cacheOut_r_valid_i & 2'h2 == sramSel; // @[Cache.scala 341:102]
  wire  _io_SRAMIO_3_cen_T_4 = isMiss & io_cacheOut_r_valid_i & 2'h3 == sramSel; // @[Cache.scala 341:102]
  assign io_cacheOut_ar_valid_o = cacheState == 2'h1; // @[Cache.scala 215:27]
  assign io_cacheOut_ar_addr_o = {io_cacheOut_ar_addr_o_hi,4'h0}; // @[Cat.scala 30:58]
  assign io_cacheOut_ar_len_o = {{7'd0}, isMiss}; // @[Cache.scala 215:27]
  assign io_cacheOut_w_valid_o = _IdleMux_T_1 & io_cacheIn_wen & isIdle; // @[Cache.scala 331:77]
  assign io_cacheOut_w_data_o = io_cacheIn_data_write; // @[Cache.scala 332:24]
  assign io_cacheOut_w_addr_o = io_cacheIn_addr; // @[Cache.scala 333:24]
  assign io_cacheOut_w_mask_o = io_cacheIn_mask; // @[Cache.scala 334:24]
  assign io_cacheOut_wsize = io_cacheIn_rsize; // @[Cache.scala 359:21]
  assign io_cacheIn_ready = isWrite & io_cacheOut_w_ready_i | isBlock | isIdle & hit & ~io_cacheIn_wen; // @[Cache.scala 357:67]
  assign io_cacheIn_data_read = offset[3] ? waysel[127:64] : waysel[63:0]; // @[Cache.scala 263:30]
  assign io_SRAMIO_0_cen = ~(io_cacheIn_valid & hitArray_0 & isIdle | isMiss & io_cacheOut_r_valid_i & 2'h0 == sramSel); // @[Cache.scala 341:16]
  assign io_SRAMIO_0_wen = ~(io_cacheIn_wen & isIdle | _io_SRAMIO_0_cen_T_4); // @[Cache.scala 343:16]
  assign io_SRAMIO_0_wdata = isMiss ? _io_SRAMIO_0_wdata_T_2 : _io_SRAMIO_0_wdata_T_6; // @[Cache.scala 344:21]
  assign io_SRAMIO_0_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  assign io_SRAMIO_0_wmask = isMiss ? _io_SRAMIO_0_wmask_T_2 : ramMaskWrite; // @[Cache.scala 349:21]
  assign io_SRAMIO_1_cen = ~(io_cacheIn_valid & hitArray_1 & isIdle | isMiss & io_cacheOut_r_valid_i & 2'h1 == sramSel); // @[Cache.scala 341:16]
  assign io_SRAMIO_1_wen = ~(io_cacheIn_wen & isIdle | _io_SRAMIO_1_cen_T_4); // @[Cache.scala 343:16]
  assign io_SRAMIO_1_wdata = isMiss ? _io_SRAMIO_0_wdata_T_2 : _io_SRAMIO_0_wdata_T_6; // @[Cache.scala 344:21]
  assign io_SRAMIO_1_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  assign io_SRAMIO_1_wmask = isMiss ? _io_SRAMIO_0_wmask_T_2 : ramMaskWrite; // @[Cache.scala 349:21]
  assign io_SRAMIO_2_cen = ~(io_cacheIn_valid & hitArray_2 & isIdle | isMiss & io_cacheOut_r_valid_i & 2'h2 == sramSel); // @[Cache.scala 341:16]
  assign io_SRAMIO_2_wen = ~(io_cacheIn_wen & isIdle | _io_SRAMIO_2_cen_T_4); // @[Cache.scala 343:16]
  assign io_SRAMIO_2_wdata = isMiss ? _io_SRAMIO_0_wdata_T_2 : _io_SRAMIO_0_wdata_T_6; // @[Cache.scala 344:21]
  assign io_SRAMIO_2_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  assign io_SRAMIO_2_wmask = isMiss ? _io_SRAMIO_0_wmask_T_2 : ramMaskWrite; // @[Cache.scala 349:21]
  assign io_SRAMIO_3_cen = ~(io_cacheIn_valid & hitArray_3 & isIdle | isMiss & io_cacheOut_r_valid_i & 2'h3 == sramSel); // @[Cache.scala 341:16]
  assign io_SRAMIO_3_wen = ~(io_cacheIn_wen & isIdle | _io_SRAMIO_3_cen_T_4); // @[Cache.scala 343:16]
  assign io_SRAMIO_3_wdata = isMiss ? _io_SRAMIO_0_wdata_T_2 : _io_SRAMIO_0_wdata_T_6; // @[Cache.scala 344:21]
  assign io_SRAMIO_3_addr = io_cacheIn_addr[9:4]; // @[Cache.scala 174:30]
  assign io_SRAMIO_3_wmask = isMiss ? _io_SRAMIO_0_wmask_T_2 : ramMaskWrite; // @[Cache.scala 349:21]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 178:27]
      cacheState <= 2'h0; // @[Cache.scala 178:27]
    end else if (2'h3 == cacheState) begin // @[Mux.scala 80:57]
      cacheState <= _writeMux_T;
    end else if (2'h2 == cacheState) begin // @[Mux.scala 80:57]
      if (io_cacheOut_w_ready_i) begin // @[Cache.scala 195:21]
        cacheState <= _writeMux_T;
      end else begin
        cacheState <= 2'h2;
      end
    end else if (2'h1 == cacheState) begin // @[Mux.scala 80:57]
      cacheState <= missMux;
    end else begin
      cacheState <= IdleMux;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_63_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_0_r <= _GEN_569;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_62_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_0_r <= _GEN_560;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_61_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_0_r <= _GEN_551;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_60_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_0_r <= _GEN_542;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_59_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_0_r <= _GEN_533;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_58_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_0_r <= _GEN_524;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_57_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_0_r <= _GEN_515;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_56_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_0_r <= _GEN_506;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_55_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_0_r <= _GEN_497;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_54_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_0_r <= _GEN_488;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_53_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_0_r <= _GEN_479;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_52_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_0_r <= _GEN_470;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_51_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_0_r <= _GEN_461;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_50_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_0_r <= _GEN_452;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_49_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_0_r <= _GEN_443;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_48_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_0_r <= _GEN_434;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_47_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_0_r <= _GEN_425;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_46_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_0_r <= _GEN_416;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_45_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_0_r <= _GEN_407;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_44_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_0_r <= _GEN_398;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_43_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_0_r <= _GEN_389;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_42_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_0_r <= _GEN_380;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_41_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_0_r <= _GEN_371;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_40_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_0_r <= _GEN_362;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_39_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_0_r <= _GEN_353;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_38_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_0_r <= _GEN_344;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_37_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_0_r <= _GEN_335;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_36_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_0_r <= _GEN_326;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_35_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_0_r <= _GEN_317;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_34_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_0_r <= _GEN_308;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_33_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_0_r <= _GEN_299;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_32_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_0_r <= _GEN_290;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_31_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_0_r <= _GEN_281;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_30_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_0_r <= _GEN_272;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_29_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_0_r <= _GEN_263;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_28_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_0_r <= _GEN_254;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_27_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_0_r <= _GEN_245;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_26_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_0_r <= _GEN_236;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_25_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_0_r <= _GEN_227;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_24_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_0_r <= _GEN_218;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_23_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_0_r <= _GEN_209;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_22_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_0_r <= _GEN_200;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_21_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_0_r <= _GEN_191;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_20_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_0_r <= _GEN_182;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_19_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_0_r <= _GEN_173;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_18_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_0_r <= _GEN_164;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_17_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_0_r <= _GEN_155;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_16_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_0_r <= _GEN_146;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_15_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_0_r <= _GEN_137;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_14_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_0_r <= _GEN_128;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_13_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_0_r <= _GEN_119;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_12_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_0_r <= _GEN_110;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_11_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_0_r <= _GEN_101;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_10_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_0_r <= _GEN_92;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_9_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_0_r <= _GEN_83;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_8_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_0_r <= _GEN_74;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_7_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_0_r <= _GEN_65;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_6_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_0_r <= _GEN_56;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_5_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_0_r <= _GEN_47;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_4_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_0_r <= _GEN_38;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_3_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_0_r <= _GEN_29;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_2_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_0_r <= _GEN_20;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_1_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_0_r <= _GEN_11;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_0_0_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_0_r <= _GEN_2;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_0_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_0_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_0_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_63_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_1_r <= _GEN_571;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_62_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_1_r <= _GEN_562;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_61_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_1_r <= _GEN_553;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_60_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_1_r <= _GEN_544;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_59_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_1_r <= _GEN_535;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_58_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_1_r <= _GEN_526;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_57_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_1_r <= _GEN_517;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_56_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_1_r <= _GEN_508;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_55_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_1_r <= _GEN_499;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_54_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_1_r <= _GEN_490;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_53_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_1_r <= _GEN_481;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_52_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_1_r <= _GEN_472;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_51_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_1_r <= _GEN_463;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_50_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_1_r <= _GEN_454;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_49_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_1_r <= _GEN_445;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_48_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_1_r <= _GEN_436;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_47_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_1_r <= _GEN_427;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_46_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_1_r <= _GEN_418;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_45_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_1_r <= _GEN_409;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_44_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_1_r <= _GEN_400;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_43_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_1_r <= _GEN_391;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_42_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_1_r <= _GEN_382;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_41_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_1_r <= _GEN_373;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_40_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_1_r <= _GEN_364;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_39_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_1_r <= _GEN_355;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_38_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_1_r <= _GEN_346;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_37_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_1_r <= _GEN_337;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_36_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_1_r <= _GEN_328;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_35_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_1_r <= _GEN_319;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_34_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_1_r <= _GEN_310;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_33_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_1_r <= _GEN_301;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_32_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_1_r <= _GEN_292;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_31_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_1_r <= _GEN_283;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_30_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_1_r <= _GEN_274;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_29_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_1_r <= _GEN_265;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_28_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_1_r <= _GEN_256;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_27_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_1_r <= _GEN_247;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_26_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_1_r <= _GEN_238;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_25_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_1_r <= _GEN_229;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_24_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_1_r <= _GEN_220;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_23_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_1_r <= _GEN_211;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_22_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_1_r <= _GEN_202;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_21_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_1_r <= _GEN_193;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_20_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_1_r <= _GEN_184;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_19_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_1_r <= _GEN_175;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_18_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_1_r <= _GEN_166;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_17_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_1_r <= _GEN_157;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_16_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_1_r <= _GEN_148;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_15_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_1_r <= _GEN_139;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_14_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_1_r <= _GEN_130;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_13_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_1_r <= _GEN_121;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_12_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_1_r <= _GEN_112;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_11_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_1_r <= _GEN_103;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_10_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_1_r <= _GEN_94;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_9_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_1_r <= _GEN_85;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_8_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_1_r <= _GEN_76;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_7_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_1_r <= _GEN_67;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_6_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_1_r <= _GEN_58;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_5_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_1_r <= _GEN_49;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_4_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_1_r <= _GEN_40;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_3_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_1_r <= _GEN_31;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_2_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_1_r <= _GEN_22;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_1_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_1_r <= _GEN_13;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_0_1_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_1_r <= _GEN_4;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_1_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_1_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_1_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_63_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_2_r <= _GEN_573;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_62_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_2_r <= _GEN_564;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_61_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_2_r <= _GEN_555;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_60_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_2_r <= _GEN_546;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_59_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_2_r <= _GEN_537;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_58_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_2_r <= _GEN_528;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_57_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_2_r <= _GEN_519;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_56_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_2_r <= _GEN_510;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_55_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_2_r <= _GEN_501;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_54_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_2_r <= _GEN_492;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_53_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_2_r <= _GEN_483;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_52_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_2_r <= _GEN_474;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_51_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_2_r <= _GEN_465;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_50_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_2_r <= _GEN_456;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_49_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_2_r <= _GEN_447;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_48_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_2_r <= _GEN_438;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_47_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_2_r <= _GEN_429;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_46_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_2_r <= _GEN_420;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_45_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_2_r <= _GEN_411;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_44_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_2_r <= _GEN_402;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_43_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_2_r <= _GEN_393;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_42_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_2_r <= _GEN_384;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_41_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_2_r <= _GEN_375;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_40_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_2_r <= _GEN_366;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_39_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_2_r <= _GEN_357;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_38_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_2_r <= _GEN_348;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_37_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_2_r <= _GEN_339;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_36_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_2_r <= _GEN_330;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_35_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_2_r <= _GEN_321;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_34_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_2_r <= _GEN_312;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_33_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_2_r <= _GEN_303;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_32_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_2_r <= _GEN_294;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_31_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_2_r <= _GEN_285;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_30_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_2_r <= _GEN_276;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_29_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_2_r <= _GEN_267;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_28_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_2_r <= _GEN_258;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_27_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_2_r <= _GEN_249;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_26_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_2_r <= _GEN_240;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_25_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_2_r <= _GEN_231;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_24_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_2_r <= _GEN_222;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_23_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_2_r <= _GEN_213;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_22_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_2_r <= _GEN_204;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_21_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_2_r <= _GEN_195;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_20_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_2_r <= _GEN_186;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_19_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_2_r <= _GEN_177;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_18_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_2_r <= _GEN_168;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_17_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_2_r <= _GEN_159;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_16_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_2_r <= _GEN_150;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_15_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_2_r <= _GEN_141;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_14_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_2_r <= _GEN_132;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_13_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_2_r <= _GEN_123;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_12_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_2_r <= _GEN_114;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_11_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_2_r <= _GEN_105;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_10_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_2_r <= _GEN_96;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_9_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_2_r <= _GEN_87;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_8_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_2_r <= _GEN_78;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_7_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_2_r <= _GEN_69;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_6_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_2_r <= _GEN_60;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_5_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_2_r <= _GEN_51;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_4_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_2_r <= _GEN_42;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_3_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_2_r <= _GEN_33;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_2_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_2_r <= _GEN_24;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_1_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_2_r <= _GEN_15;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_0_2_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_2_r <= _GEN_6;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_2_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_2_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_2_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_63_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_63_3_r <= _GEN_575;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_62_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_62_3_r <= _GEN_566;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_61_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_61_3_r <= _GEN_557;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_60_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_60_3_r <= _GEN_548;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_59_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_59_3_r <= _GEN_539;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_58_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_58_3_r <= _GEN_530;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_57_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_57_3_r <= _GEN_521;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_56_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_56_3_r <= _GEN_512;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_55_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_55_3_r <= _GEN_503;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_54_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_54_3_r <= _GEN_494;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_53_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_53_3_r <= _GEN_485;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_52_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_52_3_r <= _GEN_476;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_51_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_51_3_r <= _GEN_467;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_50_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_50_3_r <= _GEN_458;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_49_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_49_3_r <= _GEN_449;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_48_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_48_3_r <= _GEN_440;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_47_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_47_3_r <= _GEN_431;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_46_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_46_3_r <= _GEN_422;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_45_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_45_3_r <= _GEN_413;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_44_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_44_3_r <= _GEN_404;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_43_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_43_3_r <= _GEN_395;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_42_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_42_3_r <= _GEN_386;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_41_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_41_3_r <= _GEN_377;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_40_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_40_3_r <= _GEN_368;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_39_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_39_3_r <= _GEN_359;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_38_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_38_3_r <= _GEN_350;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_37_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_37_3_r <= _GEN_341;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_36_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_36_3_r <= _GEN_332;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_35_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_35_3_r <= _GEN_323;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_34_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_34_3_r <= _GEN_314;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_33_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_33_3_r <= _GEN_305;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_32_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_32_3_r <= _GEN_296;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_31_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_31_3_r <= _GEN_287;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_30_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_30_3_r <= _GEN_278;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_29_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_29_3_r <= _GEN_269;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_28_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_28_3_r <= _GEN_260;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_27_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_27_3_r <= _GEN_251;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_26_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_26_3_r <= _GEN_242;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_25_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_25_3_r <= _GEN_233;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_24_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_24_3_r <= _GEN_224;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_23_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_23_3_r <= _GEN_215;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_22_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_22_3_r <= _GEN_206;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_21_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_21_3_r <= _GEN_197;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_20_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_20_3_r <= _GEN_188;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_19_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_19_3_r <= _GEN_179;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_18_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_18_3_r <= _GEN_170;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_17_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_17_3_r <= _GEN_161;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_16_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_16_3_r <= _GEN_152;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_15_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_15_3_r <= _GEN_143;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_14_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_14_3_r <= _GEN_134;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_13_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_13_3_r <= _GEN_125;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_12_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_12_3_r <= _GEN_116;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_11_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_11_3_r <= _GEN_107;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_10_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_10_3_r <= _GEN_98;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_9_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_9_3_r <= _GEN_89;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_8_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_8_3_r <= _GEN_80;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_7_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_7_3_r <= _GEN_71;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_6_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_6_3_r <= _GEN_62;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_5_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_5_3_r <= _GEN_53;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_4_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_4_3_r <= _GEN_44;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_3_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_3_3_r <= _GEN_35;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_2_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_2_3_r <= _GEN_26;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_1_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_1_3_r <= _GEN_17;
    end
    if (reset) begin // @[Reg.scala 27:20]
      vArrayWire_0_3_r <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      vArrayWire_0_3_r <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_63_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_63_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_63_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_62_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_62_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_62_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_61_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_61_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_61_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_60_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_60_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_60_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_59_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_59_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_59_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_58_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_58_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_58_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_57_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_57_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_57_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_56_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_56_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_56_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_55_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_55_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_55_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_54_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_54_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_54_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_53_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_53_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_53_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_52_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_52_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_52_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_51_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_51_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_51_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_50_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_50_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_50_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_49_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_49_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_49_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_48_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_48_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_48_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_47_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_47_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_47_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_46_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_46_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_46_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_45_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_45_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_45_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_44_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_44_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_44_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_43_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_43_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_43_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_42_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_42_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_42_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_41_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_41_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_41_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_40_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_40_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_40_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_39_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_39_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_39_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_38_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_38_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_38_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_37_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_37_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_37_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_36_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_36_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_36_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_35_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_35_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_35_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_34_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_34_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_34_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_33_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_33_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_33_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_32_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_32_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_32_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_31_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_31_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_31_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_30_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_30_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_30_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_29_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_29_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_29_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_28_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_28_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_28_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_27_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_27_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_27_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_26_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_26_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_26_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_25_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_25_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_25_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_24_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_24_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_24_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_23_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_23_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_23_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_22_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_22_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_22_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_21_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_21_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_21_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_20_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_20_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_20_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_19_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_19_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_19_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_18_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_18_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_18_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_17_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_17_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_17_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_16_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_16_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_16_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_15_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_15_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_15_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_14_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_14_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_14_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_13_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_13_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_13_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_12_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_12_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_12_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_11_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_11_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_11_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_10_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_10_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_10_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_9_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_9_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_9_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_8_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_8_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_8_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_7_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_7_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_7_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_6_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_6_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_6_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_5_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_5_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_5_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_4_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_4_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_4_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_3_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_3_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_3_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_2_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_2_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_2_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_1_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_1_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_1_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      tagArrayWire_0_3_r <= 22'h0; // @[Reg.scala 27:20]
    end else if (_tagArrayWire_0_3_T_4) begin // @[Reg.scala 28:19]
      tagArrayWire_0_3_r <= tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_1_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_1_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_1_r <= _selArrayWire_1_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_0_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_0_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_0_r <= _selArrayWire_0_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_2_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_2_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_2_r <= _selArrayWire_2_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_3_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_3_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_3_r <= _selArrayWire_3_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_4_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_4_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_4_r <= _selArrayWire_4_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_5_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_5_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_5_r <= _selArrayWire_5_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_6_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_6_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_6_r <= _selArrayWire_6_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_7_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_7_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_7_r <= _selArrayWire_7_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_8_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_8_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_8_r <= _selArrayWire_8_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_9_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_9_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_9_r <= _selArrayWire_9_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_10_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_10_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_10_r <= _selArrayWire_10_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_11_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_11_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_11_r <= _selArrayWire_11_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_12_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_12_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_12_r <= _selArrayWire_12_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_13_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_13_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_13_r <= _selArrayWire_13_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_14_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_14_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_14_r <= _selArrayWire_14_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_15_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_15_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_15_r <= _selArrayWire_15_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_16_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_16_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_16_r <= _selArrayWire_16_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_17_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_17_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_17_r <= _selArrayWire_17_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_18_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_18_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_18_r <= _selArrayWire_18_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_19_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_19_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_19_r <= _selArrayWire_19_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_20_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_20_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_20_r <= _selArrayWire_20_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_21_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_21_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_21_r <= _selArrayWire_21_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_22_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_22_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_22_r <= _selArrayWire_22_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_23_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_23_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_23_r <= _selArrayWire_23_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_24_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_24_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_24_r <= _selArrayWire_24_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_25_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_25_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_25_r <= _selArrayWire_25_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_26_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_26_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_26_r <= _selArrayWire_26_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_27_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_27_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_27_r <= _selArrayWire_27_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_28_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_28_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_28_r <= _selArrayWire_28_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_29_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_29_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_29_r <= _selArrayWire_29_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_30_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_30_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_30_r <= _selArrayWire_30_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_31_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_31_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_31_r <= _selArrayWire_31_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_32_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_32_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_32_r <= _selArrayWire_32_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_33_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_33_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_33_r <= _selArrayWire_33_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_34_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_34_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_34_r <= _selArrayWire_34_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_35_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_35_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_35_r <= _selArrayWire_35_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_36_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_36_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_36_r <= _selArrayWire_36_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_37_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_37_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_37_r <= _selArrayWire_37_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_38_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_38_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_38_r <= _selArrayWire_38_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_39_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_39_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_39_r <= _selArrayWire_39_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_40_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_40_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_40_r <= _selArrayWire_40_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_41_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_41_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_41_r <= _selArrayWire_41_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_42_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_42_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_42_r <= _selArrayWire_42_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_43_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_43_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_43_r <= _selArrayWire_43_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_44_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_44_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_44_r <= _selArrayWire_44_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_45_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_45_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_45_r <= _selArrayWire_45_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_46_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_46_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_46_r <= _selArrayWire_46_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_47_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_47_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_47_r <= _selArrayWire_47_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_48_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_48_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_48_r <= _selArrayWire_48_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_49_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_49_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_49_r <= _selArrayWire_49_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_50_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_50_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_50_r <= _selArrayWire_50_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_51_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_51_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_51_r <= _selArrayWire_51_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_52_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_52_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_52_r <= _selArrayWire_52_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_53_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_53_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_53_r <= _selArrayWire_53_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_54_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_54_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_54_r <= _selArrayWire_54_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_55_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_55_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_55_r <= _selArrayWire_55_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_56_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_56_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_56_r <= _selArrayWire_56_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_57_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_57_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_57_r <= _selArrayWire_57_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_58_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_58_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_58_r <= _selArrayWire_58_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_59_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_59_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_59_r <= _selArrayWire_59_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_60_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_60_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_60_r <= _selArrayWire_60_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_61_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_61_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_61_r <= _selArrayWire_61_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_62_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_62_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_62_r <= _selArrayWire_62_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      selArrayWire_63_r <= 2'h0; // @[Reg.scala 27:20]
    end else if (_selArrayWire_63_T_3) begin // @[Reg.scala 28:19]
      selArrayWire_63_r <= _selArrayWire_63_T_1; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cacheState = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  vArrayWire_63_0_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vArrayWire_62_0_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  vArrayWire_61_0_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  vArrayWire_60_0_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vArrayWire_59_0_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  vArrayWire_58_0_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  vArrayWire_57_0_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  vArrayWire_56_0_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  vArrayWire_55_0_r = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  vArrayWire_54_0_r = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vArrayWire_53_0_r = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  vArrayWire_52_0_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  vArrayWire_51_0_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  vArrayWire_50_0_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  vArrayWire_49_0_r = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  vArrayWire_48_0_r = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  vArrayWire_47_0_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  vArrayWire_46_0_r = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  vArrayWire_45_0_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  vArrayWire_44_0_r = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  vArrayWire_43_0_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  vArrayWire_42_0_r = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  vArrayWire_41_0_r = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  vArrayWire_40_0_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  vArrayWire_39_0_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  vArrayWire_38_0_r = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vArrayWire_37_0_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  vArrayWire_36_0_r = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  vArrayWire_35_0_r = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  vArrayWire_34_0_r = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  vArrayWire_33_0_r = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  vArrayWire_32_0_r = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  vArrayWire_31_0_r = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  vArrayWire_30_0_r = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  vArrayWire_29_0_r = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  vArrayWire_28_0_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  vArrayWire_27_0_r = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  vArrayWire_26_0_r = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  vArrayWire_25_0_r = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  vArrayWire_24_0_r = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  vArrayWire_23_0_r = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  vArrayWire_22_0_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  vArrayWire_21_0_r = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  vArrayWire_20_0_r = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  vArrayWire_19_0_r = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  vArrayWire_18_0_r = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  vArrayWire_17_0_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  vArrayWire_16_0_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  vArrayWire_15_0_r = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  vArrayWire_14_0_r = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  vArrayWire_13_0_r = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  vArrayWire_12_0_r = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vArrayWire_11_0_r = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  vArrayWire_10_0_r = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  vArrayWire_9_0_r = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  vArrayWire_8_0_r = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  vArrayWire_7_0_r = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  vArrayWire_6_0_r = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  vArrayWire_5_0_r = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  vArrayWire_4_0_r = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  vArrayWire_3_0_r = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  vArrayWire_2_0_r = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  vArrayWire_1_0_r = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  vArrayWire_0_0_r = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tagArrayWire_63_0_r = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tagArrayWire_62_0_r = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tagArrayWire_61_0_r = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tagArrayWire_60_0_r = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tagArrayWire_59_0_r = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tagArrayWire_58_0_r = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tagArrayWire_57_0_r = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tagArrayWire_56_0_r = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tagArrayWire_55_0_r = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tagArrayWire_54_0_r = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tagArrayWire_53_0_r = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tagArrayWire_52_0_r = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tagArrayWire_51_0_r = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tagArrayWire_50_0_r = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tagArrayWire_49_0_r = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tagArrayWire_48_0_r = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tagArrayWire_47_0_r = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tagArrayWire_46_0_r = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tagArrayWire_45_0_r = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tagArrayWire_44_0_r = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tagArrayWire_43_0_r = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tagArrayWire_42_0_r = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tagArrayWire_41_0_r = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tagArrayWire_40_0_r = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tagArrayWire_39_0_r = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tagArrayWire_38_0_r = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tagArrayWire_37_0_r = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tagArrayWire_36_0_r = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tagArrayWire_35_0_r = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tagArrayWire_34_0_r = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tagArrayWire_33_0_r = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tagArrayWire_32_0_r = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tagArrayWire_31_0_r = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tagArrayWire_30_0_r = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tagArrayWire_29_0_r = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tagArrayWire_28_0_r = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tagArrayWire_27_0_r = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tagArrayWire_26_0_r = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tagArrayWire_25_0_r = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tagArrayWire_24_0_r = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tagArrayWire_23_0_r = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tagArrayWire_22_0_r = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tagArrayWire_21_0_r = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tagArrayWire_20_0_r = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tagArrayWire_19_0_r = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tagArrayWire_18_0_r = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tagArrayWire_17_0_r = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tagArrayWire_16_0_r = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tagArrayWire_15_0_r = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tagArrayWire_14_0_r = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tagArrayWire_13_0_r = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tagArrayWire_12_0_r = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tagArrayWire_11_0_r = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tagArrayWire_10_0_r = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tagArrayWire_9_0_r = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tagArrayWire_8_0_r = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tagArrayWire_7_0_r = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tagArrayWire_6_0_r = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tagArrayWire_5_0_r = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tagArrayWire_4_0_r = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tagArrayWire_3_0_r = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tagArrayWire_2_0_r = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tagArrayWire_1_0_r = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  tagArrayWire_0_0_r = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  vArrayWire_63_1_r = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  vArrayWire_62_1_r = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  vArrayWire_61_1_r = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  vArrayWire_60_1_r = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  vArrayWire_59_1_r = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  vArrayWire_58_1_r = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  vArrayWire_57_1_r = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  vArrayWire_56_1_r = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  vArrayWire_55_1_r = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  vArrayWire_54_1_r = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  vArrayWire_53_1_r = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  vArrayWire_52_1_r = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  vArrayWire_51_1_r = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  vArrayWire_50_1_r = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  vArrayWire_49_1_r = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  vArrayWire_48_1_r = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  vArrayWire_47_1_r = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  vArrayWire_46_1_r = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  vArrayWire_45_1_r = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  vArrayWire_44_1_r = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  vArrayWire_43_1_r = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  vArrayWire_42_1_r = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  vArrayWire_41_1_r = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  vArrayWire_40_1_r = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  vArrayWire_39_1_r = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  vArrayWire_38_1_r = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  vArrayWire_37_1_r = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  vArrayWire_36_1_r = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  vArrayWire_35_1_r = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  vArrayWire_34_1_r = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  vArrayWire_33_1_r = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  vArrayWire_32_1_r = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  vArrayWire_31_1_r = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  vArrayWire_30_1_r = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  vArrayWire_29_1_r = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  vArrayWire_28_1_r = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  vArrayWire_27_1_r = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  vArrayWire_26_1_r = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  vArrayWire_25_1_r = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  vArrayWire_24_1_r = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  vArrayWire_23_1_r = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  vArrayWire_22_1_r = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  vArrayWire_21_1_r = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  vArrayWire_20_1_r = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  vArrayWire_19_1_r = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  vArrayWire_18_1_r = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  vArrayWire_17_1_r = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  vArrayWire_16_1_r = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  vArrayWire_15_1_r = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  vArrayWire_14_1_r = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  vArrayWire_13_1_r = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  vArrayWire_12_1_r = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  vArrayWire_11_1_r = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  vArrayWire_10_1_r = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vArrayWire_9_1_r = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  vArrayWire_8_1_r = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  vArrayWire_7_1_r = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  vArrayWire_6_1_r = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  vArrayWire_5_1_r = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  vArrayWire_4_1_r = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  vArrayWire_3_1_r = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  vArrayWire_2_1_r = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  vArrayWire_1_1_r = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  vArrayWire_0_1_r = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tagArrayWire_63_1_r = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  tagArrayWire_62_1_r = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  tagArrayWire_61_1_r = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  tagArrayWire_60_1_r = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  tagArrayWire_59_1_r = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  tagArrayWire_58_1_r = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  tagArrayWire_57_1_r = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  tagArrayWire_56_1_r = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  tagArrayWire_55_1_r = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  tagArrayWire_54_1_r = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  tagArrayWire_53_1_r = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  tagArrayWire_52_1_r = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  tagArrayWire_51_1_r = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  tagArrayWire_50_1_r = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  tagArrayWire_49_1_r = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  tagArrayWire_48_1_r = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  tagArrayWire_47_1_r = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  tagArrayWire_46_1_r = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  tagArrayWire_45_1_r = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  tagArrayWire_44_1_r = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  tagArrayWire_43_1_r = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  tagArrayWire_42_1_r = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  tagArrayWire_41_1_r = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  tagArrayWire_40_1_r = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  tagArrayWire_39_1_r = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  tagArrayWire_38_1_r = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  tagArrayWire_37_1_r = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  tagArrayWire_36_1_r = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  tagArrayWire_35_1_r = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  tagArrayWire_34_1_r = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  tagArrayWire_33_1_r = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  tagArrayWire_32_1_r = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  tagArrayWire_31_1_r = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  tagArrayWire_30_1_r = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  tagArrayWire_29_1_r = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  tagArrayWire_28_1_r = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  tagArrayWire_27_1_r = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  tagArrayWire_26_1_r = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  tagArrayWire_25_1_r = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  tagArrayWire_24_1_r = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  tagArrayWire_23_1_r = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  tagArrayWire_22_1_r = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  tagArrayWire_21_1_r = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  tagArrayWire_20_1_r = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  tagArrayWire_19_1_r = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  tagArrayWire_18_1_r = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  tagArrayWire_17_1_r = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  tagArrayWire_16_1_r = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  tagArrayWire_15_1_r = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  tagArrayWire_14_1_r = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  tagArrayWire_13_1_r = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  tagArrayWire_12_1_r = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  tagArrayWire_11_1_r = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  tagArrayWire_10_1_r = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  tagArrayWire_9_1_r = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  tagArrayWire_8_1_r = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  tagArrayWire_7_1_r = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  tagArrayWire_6_1_r = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  tagArrayWire_5_1_r = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  tagArrayWire_4_1_r = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  tagArrayWire_3_1_r = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  tagArrayWire_2_1_r = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  tagArrayWire_1_1_r = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  tagArrayWire_0_1_r = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  vArrayWire_63_2_r = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  vArrayWire_62_2_r = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  vArrayWire_61_2_r = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  vArrayWire_60_2_r = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  vArrayWire_59_2_r = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  vArrayWire_58_2_r = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  vArrayWire_57_2_r = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  vArrayWire_56_2_r = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  vArrayWire_55_2_r = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  vArrayWire_54_2_r = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  vArrayWire_53_2_r = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  vArrayWire_52_2_r = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  vArrayWire_51_2_r = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  vArrayWire_50_2_r = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  vArrayWire_49_2_r = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  vArrayWire_48_2_r = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  vArrayWire_47_2_r = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  vArrayWire_46_2_r = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  vArrayWire_45_2_r = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  vArrayWire_44_2_r = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  vArrayWire_43_2_r = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  vArrayWire_42_2_r = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  vArrayWire_41_2_r = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  vArrayWire_40_2_r = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  vArrayWire_39_2_r = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  vArrayWire_38_2_r = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  vArrayWire_37_2_r = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  vArrayWire_36_2_r = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  vArrayWire_35_2_r = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  vArrayWire_34_2_r = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  vArrayWire_33_2_r = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  vArrayWire_32_2_r = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  vArrayWire_31_2_r = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  vArrayWire_30_2_r = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  vArrayWire_29_2_r = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  vArrayWire_28_2_r = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  vArrayWire_27_2_r = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  vArrayWire_26_2_r = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  vArrayWire_25_2_r = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  vArrayWire_24_2_r = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  vArrayWire_23_2_r = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  vArrayWire_22_2_r = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  vArrayWire_21_2_r = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  vArrayWire_20_2_r = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  vArrayWire_19_2_r = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  vArrayWire_18_2_r = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  vArrayWire_17_2_r = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  vArrayWire_16_2_r = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  vArrayWire_15_2_r = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  vArrayWire_14_2_r = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  vArrayWire_13_2_r = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  vArrayWire_12_2_r = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  vArrayWire_11_2_r = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  vArrayWire_10_2_r = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  vArrayWire_9_2_r = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  vArrayWire_8_2_r = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  vArrayWire_7_2_r = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  vArrayWire_6_2_r = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  vArrayWire_5_2_r = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  vArrayWire_4_2_r = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  vArrayWire_3_2_r = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  vArrayWire_2_2_r = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  vArrayWire_1_2_r = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  vArrayWire_0_2_r = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  tagArrayWire_63_2_r = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  tagArrayWire_62_2_r = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  tagArrayWire_61_2_r = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  tagArrayWire_60_2_r = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  tagArrayWire_59_2_r = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  tagArrayWire_58_2_r = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  tagArrayWire_57_2_r = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  tagArrayWire_56_2_r = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  tagArrayWire_55_2_r = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  tagArrayWire_54_2_r = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  tagArrayWire_53_2_r = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  tagArrayWire_52_2_r = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  tagArrayWire_51_2_r = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  tagArrayWire_50_2_r = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  tagArrayWire_49_2_r = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  tagArrayWire_48_2_r = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  tagArrayWire_47_2_r = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  tagArrayWire_46_2_r = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  tagArrayWire_45_2_r = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  tagArrayWire_44_2_r = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  tagArrayWire_43_2_r = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  tagArrayWire_42_2_r = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  tagArrayWire_41_2_r = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  tagArrayWire_40_2_r = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  tagArrayWire_39_2_r = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  tagArrayWire_38_2_r = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  tagArrayWire_37_2_r = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  tagArrayWire_36_2_r = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  tagArrayWire_35_2_r = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  tagArrayWire_34_2_r = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  tagArrayWire_33_2_r = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  tagArrayWire_32_2_r = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  tagArrayWire_31_2_r = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  tagArrayWire_30_2_r = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  tagArrayWire_29_2_r = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  tagArrayWire_28_2_r = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  tagArrayWire_27_2_r = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  tagArrayWire_26_2_r = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  tagArrayWire_25_2_r = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  tagArrayWire_24_2_r = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  tagArrayWire_23_2_r = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  tagArrayWire_22_2_r = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  tagArrayWire_21_2_r = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  tagArrayWire_20_2_r = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  tagArrayWire_19_2_r = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  tagArrayWire_18_2_r = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  tagArrayWire_17_2_r = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  tagArrayWire_16_2_r = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  tagArrayWire_15_2_r = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  tagArrayWire_14_2_r = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  tagArrayWire_13_2_r = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  tagArrayWire_12_2_r = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  tagArrayWire_11_2_r = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  tagArrayWire_10_2_r = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  tagArrayWire_9_2_r = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  tagArrayWire_8_2_r = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  tagArrayWire_7_2_r = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  tagArrayWire_6_2_r = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  tagArrayWire_5_2_r = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  tagArrayWire_4_2_r = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  tagArrayWire_3_2_r = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  tagArrayWire_2_2_r = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  tagArrayWire_1_2_r = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  tagArrayWire_0_2_r = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  vArrayWire_63_3_r = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  vArrayWire_62_3_r = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  vArrayWire_61_3_r = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  vArrayWire_60_3_r = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  vArrayWire_59_3_r = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  vArrayWire_58_3_r = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  vArrayWire_57_3_r = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  vArrayWire_56_3_r = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  vArrayWire_55_3_r = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  vArrayWire_54_3_r = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  vArrayWire_53_3_r = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  vArrayWire_52_3_r = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  vArrayWire_51_3_r = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  vArrayWire_50_3_r = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  vArrayWire_49_3_r = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  vArrayWire_48_3_r = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  vArrayWire_47_3_r = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  vArrayWire_46_3_r = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  vArrayWire_45_3_r = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  vArrayWire_44_3_r = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  vArrayWire_43_3_r = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  vArrayWire_42_3_r = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  vArrayWire_41_3_r = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  vArrayWire_40_3_r = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  vArrayWire_39_3_r = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  vArrayWire_38_3_r = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  vArrayWire_37_3_r = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  vArrayWire_36_3_r = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  vArrayWire_35_3_r = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  vArrayWire_34_3_r = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  vArrayWire_33_3_r = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  vArrayWire_32_3_r = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  vArrayWire_31_3_r = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  vArrayWire_30_3_r = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  vArrayWire_29_3_r = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  vArrayWire_28_3_r = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  vArrayWire_27_3_r = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  vArrayWire_26_3_r = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  vArrayWire_25_3_r = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  vArrayWire_24_3_r = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  vArrayWire_23_3_r = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  vArrayWire_22_3_r = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  vArrayWire_21_3_r = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  vArrayWire_20_3_r = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  vArrayWire_19_3_r = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  vArrayWire_18_3_r = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  vArrayWire_17_3_r = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  vArrayWire_16_3_r = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  vArrayWire_15_3_r = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  vArrayWire_14_3_r = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  vArrayWire_13_3_r = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  vArrayWire_12_3_r = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  vArrayWire_11_3_r = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  vArrayWire_10_3_r = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  vArrayWire_9_3_r = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  vArrayWire_8_3_r = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  vArrayWire_7_3_r = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  vArrayWire_6_3_r = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  vArrayWire_5_3_r = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  vArrayWire_4_3_r = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  vArrayWire_3_3_r = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  vArrayWire_2_3_r = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  vArrayWire_1_3_r = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  vArrayWire_0_3_r = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  tagArrayWire_63_3_r = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  tagArrayWire_62_3_r = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  tagArrayWire_61_3_r = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  tagArrayWire_60_3_r = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  tagArrayWire_59_3_r = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  tagArrayWire_58_3_r = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  tagArrayWire_57_3_r = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  tagArrayWire_56_3_r = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  tagArrayWire_55_3_r = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  tagArrayWire_54_3_r = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  tagArrayWire_53_3_r = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  tagArrayWire_52_3_r = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  tagArrayWire_51_3_r = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  tagArrayWire_50_3_r = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  tagArrayWire_49_3_r = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  tagArrayWire_48_3_r = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  tagArrayWire_47_3_r = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  tagArrayWire_46_3_r = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  tagArrayWire_45_3_r = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  tagArrayWire_44_3_r = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  tagArrayWire_43_3_r = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  tagArrayWire_42_3_r = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  tagArrayWire_41_3_r = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  tagArrayWire_40_3_r = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  tagArrayWire_39_3_r = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  tagArrayWire_38_3_r = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  tagArrayWire_37_3_r = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  tagArrayWire_36_3_r = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  tagArrayWire_35_3_r = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  tagArrayWire_34_3_r = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  tagArrayWire_33_3_r = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  tagArrayWire_32_3_r = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  tagArrayWire_31_3_r = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  tagArrayWire_30_3_r = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  tagArrayWire_29_3_r = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  tagArrayWire_28_3_r = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  tagArrayWire_27_3_r = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  tagArrayWire_26_3_r = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  tagArrayWire_25_3_r = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  tagArrayWire_24_3_r = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  tagArrayWire_23_3_r = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  tagArrayWire_22_3_r = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  tagArrayWire_21_3_r = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  tagArrayWire_20_3_r = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  tagArrayWire_19_3_r = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  tagArrayWire_18_3_r = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  tagArrayWire_17_3_r = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  tagArrayWire_16_3_r = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  tagArrayWire_15_3_r = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  tagArrayWire_14_3_r = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  tagArrayWire_13_3_r = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  tagArrayWire_12_3_r = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  tagArrayWire_11_3_r = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  tagArrayWire_10_3_r = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  tagArrayWire_9_3_r = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  tagArrayWire_8_3_r = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  tagArrayWire_7_3_r = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  tagArrayWire_6_3_r = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  tagArrayWire_5_3_r = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  tagArrayWire_4_3_r = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  tagArrayWire_3_3_r = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  tagArrayWire_2_3_r = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  tagArrayWire_1_3_r = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  tagArrayWire_0_3_r = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  selArrayWire_1_r = _RAND_513[1:0];
  _RAND_514 = {1{`RANDOM}};
  selArrayWire_0_r = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  selArrayWire_2_r = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  selArrayWire_3_r = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  selArrayWire_4_r = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  selArrayWire_5_r = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  selArrayWire_6_r = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  selArrayWire_7_r = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  selArrayWire_8_r = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  selArrayWire_9_r = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  selArrayWire_10_r = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  selArrayWire_11_r = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  selArrayWire_12_r = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  selArrayWire_13_r = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  selArrayWire_14_r = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  selArrayWire_15_r = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  selArrayWire_16_r = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  selArrayWire_17_r = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  selArrayWire_18_r = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  selArrayWire_19_r = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  selArrayWire_20_r = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  selArrayWire_21_r = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  selArrayWire_22_r = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  selArrayWire_23_r = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  selArrayWire_24_r = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  selArrayWire_25_r = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  selArrayWire_26_r = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  selArrayWire_27_r = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  selArrayWire_28_r = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  selArrayWire_29_r = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  selArrayWire_30_r = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  selArrayWire_31_r = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  selArrayWire_32_r = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  selArrayWire_33_r = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  selArrayWire_34_r = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  selArrayWire_35_r = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  selArrayWire_36_r = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  selArrayWire_37_r = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  selArrayWire_38_r = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  selArrayWire_39_r = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  selArrayWire_40_r = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  selArrayWire_41_r = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  selArrayWire_42_r = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  selArrayWire_43_r = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  selArrayWire_44_r = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  selArrayWire_45_r = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  selArrayWire_46_r = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  selArrayWire_47_r = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  selArrayWire_48_r = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  selArrayWire_49_r = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  selArrayWire_50_r = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  selArrayWire_51_r = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  selArrayWire_52_r = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  selArrayWire_53_r = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  selArrayWire_54_r = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  selArrayWire_55_r = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  selArrayWire_56_r = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  selArrayWire_57_r = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  selArrayWire_58_r = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  selArrayWire_59_r = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  selArrayWire_60_r = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  selArrayWire_61_r = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  selArrayWire_62_r = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  selArrayWire_63_r = _RAND_576[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module clint(
  input         clock,
  input         reset,
  input         io_clintIO_valid,
  output [63:0] io_clintIO_data_read,
  input  [63:0] io_clintIO_data_write,
  input         io_clintIO_wen,
  input  [31:0] io_clintIO_addr,
  output        intrTimeCnt_0,
  input         startTimeCnt_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime_r; // @[Reg.scala 27:20]
  wire [63:0] _mtime_T_1 = mtime_r + 64'h1; // @[clint.scala 21:30]
  wire  _mtimecmp_T_4 = io_clintIO_valid & io_clintIO_wen & io_clintIO_addr == 32'h2004000; // @[clint.scala 23:87]
  reg [63:0] mtimecmp_r; // @[Reg.scala 27:20]
  wire [63:0] _io_clintIO_data_read_T_5 = 32'h2004000 == io_clintIO_addr ? mtimecmp_r : 64'h0; // @[Mux.scala 80:57]
  wire  intrTimeCnt = mtime_r >= mtimecmp_r & startTimeCnt_0; // @[clint.scala 37:36]
  assign io_clintIO_data_read = 32'h200bff8 == io_clintIO_addr ? mtime_r : _io_clintIO_data_read_T_5; // @[Mux.scala 80:57]
  assign intrTimeCnt_0 = intrTimeCnt;
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      mtime_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (startTimeCnt_0) begin // @[Reg.scala 28:19]
      mtime_r <= _mtime_T_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      mtimecmp_r <= 64'h0; // @[Reg.scala 27:20]
    end else if (_mtimecmp_T_4) begin // @[Reg.scala 28:19]
      mtimecmp_r <= io_clintIO_data_write; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime_r = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp_r = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mem(
  input          clock,
  input          io_memIO_cen,
  input          io_memIO_wen,
  input  [127:0] io_memIO_wdata,
  input  [5:0]   io_memIO_addr,
  input  [127:0] io_memIO_wmask,
  output [127:0] io_memIO_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [127:0] _RAND_19;
  reg [127:0] _RAND_20;
  reg [127:0] _RAND_21;
  reg [127:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [127:0] _RAND_27;
  reg [127:0] _RAND_28;
  reg [127:0] _RAND_29;
  reg [127:0] _RAND_30;
  reg [127:0] _RAND_31;
  reg [127:0] _RAND_32;
  reg [127:0] _RAND_33;
  reg [127:0] _RAND_34;
  reg [127:0] _RAND_35;
  reg [127:0] _RAND_36;
  reg [127:0] _RAND_37;
  reg [127:0] _RAND_38;
  reg [127:0] _RAND_39;
  reg [127:0] _RAND_40;
  reg [127:0] _RAND_41;
  reg [127:0] _RAND_42;
  reg [127:0] _RAND_43;
  reg [127:0] _RAND_44;
  reg [127:0] _RAND_45;
  reg [127:0] _RAND_46;
  reg [127:0] _RAND_47;
  reg [127:0] _RAND_48;
  reg [127:0] _RAND_49;
  reg [127:0] _RAND_50;
  reg [127:0] _RAND_51;
  reg [127:0] _RAND_52;
  reg [127:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [127:0] _RAND_55;
  reg [127:0] _RAND_56;
  reg [127:0] _RAND_57;
  reg [127:0] _RAND_58;
  reg [127:0] _RAND_59;
  reg [127:0] _RAND_60;
  reg [127:0] _RAND_61;
  reg [127:0] _RAND_62;
  reg [127:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire  cen = ~io_memIO_cen; // @[mem.scala 14:14]
  wire [127:0] bwen = ~io_memIO_wmask; // @[mem.scala 15:15]
  wire  wen = ~io_memIO_wen; // @[mem.scala 16:14]
  wire [127:0] _ramWire_0_T = io_memIO_wdata & bwen; // @[mem.scala 25:47]
  reg [127:0] ramWire_0_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_0_T_1 = ramWire_0_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_0_T_2 = _ramWire_0_T | _ramWire_0_T_1; // @[mem.scala 25:55]
  wire  _ramWire_0_T_5 = cen & wen & io_memIO_addr == 6'h0; // @[mem.scala 25:98]
  reg [127:0] ramWire_1_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_1_T_1 = ramWire_1_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_1_T_2 = _ramWire_0_T | _ramWire_1_T_1; // @[mem.scala 25:55]
  wire  _ramWire_1_T_5 = cen & wen & io_memIO_addr == 6'h1; // @[mem.scala 25:98]
  reg [127:0] ramWire_2_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_2_T_1 = ramWire_2_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_2_T_2 = _ramWire_0_T | _ramWire_2_T_1; // @[mem.scala 25:55]
  wire  _ramWire_2_T_5 = cen & wen & io_memIO_addr == 6'h2; // @[mem.scala 25:98]
  reg [127:0] ramWire_3_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_3_T_1 = ramWire_3_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_3_T_2 = _ramWire_0_T | _ramWire_3_T_1; // @[mem.scala 25:55]
  wire  _ramWire_3_T_5 = cen & wen & io_memIO_addr == 6'h3; // @[mem.scala 25:98]
  reg [127:0] ramWire_4_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_4_T_1 = ramWire_4_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_4_T_2 = _ramWire_0_T | _ramWire_4_T_1; // @[mem.scala 25:55]
  wire  _ramWire_4_T_5 = cen & wen & io_memIO_addr == 6'h4; // @[mem.scala 25:98]
  reg [127:0] ramWire_5_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_5_T_1 = ramWire_5_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_5_T_2 = _ramWire_0_T | _ramWire_5_T_1; // @[mem.scala 25:55]
  wire  _ramWire_5_T_5 = cen & wen & io_memIO_addr == 6'h5; // @[mem.scala 25:98]
  reg [127:0] ramWire_6_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_6_T_1 = ramWire_6_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_6_T_2 = _ramWire_0_T | _ramWire_6_T_1; // @[mem.scala 25:55]
  wire  _ramWire_6_T_5 = cen & wen & io_memIO_addr == 6'h6; // @[mem.scala 25:98]
  reg [127:0] ramWire_7_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_7_T_1 = ramWire_7_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_7_T_2 = _ramWire_0_T | _ramWire_7_T_1; // @[mem.scala 25:55]
  wire  _ramWire_7_T_5 = cen & wen & io_memIO_addr == 6'h7; // @[mem.scala 25:98]
  reg [127:0] ramWire_8_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_8_T_1 = ramWire_8_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_8_T_2 = _ramWire_0_T | _ramWire_8_T_1; // @[mem.scala 25:55]
  wire  _ramWire_8_T_5 = cen & wen & io_memIO_addr == 6'h8; // @[mem.scala 25:98]
  reg [127:0] ramWire_9_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_9_T_1 = ramWire_9_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_9_T_2 = _ramWire_0_T | _ramWire_9_T_1; // @[mem.scala 25:55]
  wire  _ramWire_9_T_5 = cen & wen & io_memIO_addr == 6'h9; // @[mem.scala 25:98]
  reg [127:0] ramWire_10_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_10_T_1 = ramWire_10_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_10_T_2 = _ramWire_0_T | _ramWire_10_T_1; // @[mem.scala 25:55]
  wire  _ramWire_10_T_5 = cen & wen & io_memIO_addr == 6'ha; // @[mem.scala 25:98]
  reg [127:0] ramWire_11_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_11_T_1 = ramWire_11_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_11_T_2 = _ramWire_0_T | _ramWire_11_T_1; // @[mem.scala 25:55]
  wire  _ramWire_11_T_5 = cen & wen & io_memIO_addr == 6'hb; // @[mem.scala 25:98]
  reg [127:0] ramWire_12_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_12_T_1 = ramWire_12_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_12_T_2 = _ramWire_0_T | _ramWire_12_T_1; // @[mem.scala 25:55]
  wire  _ramWire_12_T_5 = cen & wen & io_memIO_addr == 6'hc; // @[mem.scala 25:98]
  reg [127:0] ramWire_13_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_13_T_1 = ramWire_13_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_13_T_2 = _ramWire_0_T | _ramWire_13_T_1; // @[mem.scala 25:55]
  wire  _ramWire_13_T_5 = cen & wen & io_memIO_addr == 6'hd; // @[mem.scala 25:98]
  reg [127:0] ramWire_14_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_14_T_1 = ramWire_14_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_14_T_2 = _ramWire_0_T | _ramWire_14_T_1; // @[mem.scala 25:55]
  wire  _ramWire_14_T_5 = cen & wen & io_memIO_addr == 6'he; // @[mem.scala 25:98]
  reg [127:0] ramWire_15_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_15_T_1 = ramWire_15_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_15_T_2 = _ramWire_0_T | _ramWire_15_T_1; // @[mem.scala 25:55]
  wire  _ramWire_15_T_5 = cen & wen & io_memIO_addr == 6'hf; // @[mem.scala 25:98]
  reg [127:0] ramWire_16_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_16_T_1 = ramWire_16_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_16_T_2 = _ramWire_0_T | _ramWire_16_T_1; // @[mem.scala 25:55]
  wire  _ramWire_16_T_5 = cen & wen & io_memIO_addr == 6'h10; // @[mem.scala 25:98]
  reg [127:0] ramWire_17_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_17_T_1 = ramWire_17_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_17_T_2 = _ramWire_0_T | _ramWire_17_T_1; // @[mem.scala 25:55]
  wire  _ramWire_17_T_5 = cen & wen & io_memIO_addr == 6'h11; // @[mem.scala 25:98]
  reg [127:0] ramWire_18_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_18_T_1 = ramWire_18_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_18_T_2 = _ramWire_0_T | _ramWire_18_T_1; // @[mem.scala 25:55]
  wire  _ramWire_18_T_5 = cen & wen & io_memIO_addr == 6'h12; // @[mem.scala 25:98]
  reg [127:0] ramWire_19_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_19_T_1 = ramWire_19_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_19_T_2 = _ramWire_0_T | _ramWire_19_T_1; // @[mem.scala 25:55]
  wire  _ramWire_19_T_5 = cen & wen & io_memIO_addr == 6'h13; // @[mem.scala 25:98]
  reg [127:0] ramWire_20_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_20_T_1 = ramWire_20_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_20_T_2 = _ramWire_0_T | _ramWire_20_T_1; // @[mem.scala 25:55]
  wire  _ramWire_20_T_5 = cen & wen & io_memIO_addr == 6'h14; // @[mem.scala 25:98]
  reg [127:0] ramWire_21_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_21_T_1 = ramWire_21_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_21_T_2 = _ramWire_0_T | _ramWire_21_T_1; // @[mem.scala 25:55]
  wire  _ramWire_21_T_5 = cen & wen & io_memIO_addr == 6'h15; // @[mem.scala 25:98]
  reg [127:0] ramWire_22_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_22_T_1 = ramWire_22_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_22_T_2 = _ramWire_0_T | _ramWire_22_T_1; // @[mem.scala 25:55]
  wire  _ramWire_22_T_5 = cen & wen & io_memIO_addr == 6'h16; // @[mem.scala 25:98]
  reg [127:0] ramWire_23_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_23_T_1 = ramWire_23_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_23_T_2 = _ramWire_0_T | _ramWire_23_T_1; // @[mem.scala 25:55]
  wire  _ramWire_23_T_5 = cen & wen & io_memIO_addr == 6'h17; // @[mem.scala 25:98]
  reg [127:0] ramWire_24_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_24_T_1 = ramWire_24_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_24_T_2 = _ramWire_0_T | _ramWire_24_T_1; // @[mem.scala 25:55]
  wire  _ramWire_24_T_5 = cen & wen & io_memIO_addr == 6'h18; // @[mem.scala 25:98]
  reg [127:0] ramWire_25_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_25_T_1 = ramWire_25_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_25_T_2 = _ramWire_0_T | _ramWire_25_T_1; // @[mem.scala 25:55]
  wire  _ramWire_25_T_5 = cen & wen & io_memIO_addr == 6'h19; // @[mem.scala 25:98]
  reg [127:0] ramWire_26_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_26_T_1 = ramWire_26_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_26_T_2 = _ramWire_0_T | _ramWire_26_T_1; // @[mem.scala 25:55]
  wire  _ramWire_26_T_5 = cen & wen & io_memIO_addr == 6'h1a; // @[mem.scala 25:98]
  reg [127:0] ramWire_27_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_27_T_1 = ramWire_27_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_27_T_2 = _ramWire_0_T | _ramWire_27_T_1; // @[mem.scala 25:55]
  wire  _ramWire_27_T_5 = cen & wen & io_memIO_addr == 6'h1b; // @[mem.scala 25:98]
  reg [127:0] ramWire_28_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_28_T_1 = ramWire_28_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_28_T_2 = _ramWire_0_T | _ramWire_28_T_1; // @[mem.scala 25:55]
  wire  _ramWire_28_T_5 = cen & wen & io_memIO_addr == 6'h1c; // @[mem.scala 25:98]
  reg [127:0] ramWire_29_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_29_T_1 = ramWire_29_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_29_T_2 = _ramWire_0_T | _ramWire_29_T_1; // @[mem.scala 25:55]
  wire  _ramWire_29_T_5 = cen & wen & io_memIO_addr == 6'h1d; // @[mem.scala 25:98]
  reg [127:0] ramWire_30_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_30_T_1 = ramWire_30_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_30_T_2 = _ramWire_0_T | _ramWire_30_T_1; // @[mem.scala 25:55]
  wire  _ramWire_30_T_5 = cen & wen & io_memIO_addr == 6'h1e; // @[mem.scala 25:98]
  reg [127:0] ramWire_31_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_31_T_1 = ramWire_31_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_31_T_2 = _ramWire_0_T | _ramWire_31_T_1; // @[mem.scala 25:55]
  wire  _ramWire_31_T_5 = cen & wen & io_memIO_addr == 6'h1f; // @[mem.scala 25:98]
  reg [127:0] ramWire_32_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_32_T_1 = ramWire_32_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_32_T_2 = _ramWire_0_T | _ramWire_32_T_1; // @[mem.scala 25:55]
  wire  _ramWire_32_T_5 = cen & wen & io_memIO_addr == 6'h20; // @[mem.scala 25:98]
  reg [127:0] ramWire_33_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_33_T_1 = ramWire_33_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_33_T_2 = _ramWire_0_T | _ramWire_33_T_1; // @[mem.scala 25:55]
  wire  _ramWire_33_T_5 = cen & wen & io_memIO_addr == 6'h21; // @[mem.scala 25:98]
  reg [127:0] ramWire_34_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_34_T_1 = ramWire_34_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_34_T_2 = _ramWire_0_T | _ramWire_34_T_1; // @[mem.scala 25:55]
  wire  _ramWire_34_T_5 = cen & wen & io_memIO_addr == 6'h22; // @[mem.scala 25:98]
  reg [127:0] ramWire_35_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_35_T_1 = ramWire_35_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_35_T_2 = _ramWire_0_T | _ramWire_35_T_1; // @[mem.scala 25:55]
  wire  _ramWire_35_T_5 = cen & wen & io_memIO_addr == 6'h23; // @[mem.scala 25:98]
  reg [127:0] ramWire_36_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_36_T_1 = ramWire_36_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_36_T_2 = _ramWire_0_T | _ramWire_36_T_1; // @[mem.scala 25:55]
  wire  _ramWire_36_T_5 = cen & wen & io_memIO_addr == 6'h24; // @[mem.scala 25:98]
  reg [127:0] ramWire_37_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_37_T_1 = ramWire_37_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_37_T_2 = _ramWire_0_T | _ramWire_37_T_1; // @[mem.scala 25:55]
  wire  _ramWire_37_T_5 = cen & wen & io_memIO_addr == 6'h25; // @[mem.scala 25:98]
  reg [127:0] ramWire_38_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_38_T_1 = ramWire_38_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_38_T_2 = _ramWire_0_T | _ramWire_38_T_1; // @[mem.scala 25:55]
  wire  _ramWire_38_T_5 = cen & wen & io_memIO_addr == 6'h26; // @[mem.scala 25:98]
  reg [127:0] ramWire_39_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_39_T_1 = ramWire_39_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_39_T_2 = _ramWire_0_T | _ramWire_39_T_1; // @[mem.scala 25:55]
  wire  _ramWire_39_T_5 = cen & wen & io_memIO_addr == 6'h27; // @[mem.scala 25:98]
  reg [127:0] ramWire_40_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_40_T_1 = ramWire_40_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_40_T_2 = _ramWire_0_T | _ramWire_40_T_1; // @[mem.scala 25:55]
  wire  _ramWire_40_T_5 = cen & wen & io_memIO_addr == 6'h28; // @[mem.scala 25:98]
  reg [127:0] ramWire_41_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_41_T_1 = ramWire_41_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_41_T_2 = _ramWire_0_T | _ramWire_41_T_1; // @[mem.scala 25:55]
  wire  _ramWire_41_T_5 = cen & wen & io_memIO_addr == 6'h29; // @[mem.scala 25:98]
  reg [127:0] ramWire_42_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_42_T_1 = ramWire_42_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_42_T_2 = _ramWire_0_T | _ramWire_42_T_1; // @[mem.scala 25:55]
  wire  _ramWire_42_T_5 = cen & wen & io_memIO_addr == 6'h2a; // @[mem.scala 25:98]
  reg [127:0] ramWire_43_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_43_T_1 = ramWire_43_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_43_T_2 = _ramWire_0_T | _ramWire_43_T_1; // @[mem.scala 25:55]
  wire  _ramWire_43_T_5 = cen & wen & io_memIO_addr == 6'h2b; // @[mem.scala 25:98]
  reg [127:0] ramWire_44_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_44_T_1 = ramWire_44_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_44_T_2 = _ramWire_0_T | _ramWire_44_T_1; // @[mem.scala 25:55]
  wire  _ramWire_44_T_5 = cen & wen & io_memIO_addr == 6'h2c; // @[mem.scala 25:98]
  reg [127:0] ramWire_45_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_45_T_1 = ramWire_45_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_45_T_2 = _ramWire_0_T | _ramWire_45_T_1; // @[mem.scala 25:55]
  wire  _ramWire_45_T_5 = cen & wen & io_memIO_addr == 6'h2d; // @[mem.scala 25:98]
  reg [127:0] ramWire_46_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_46_T_1 = ramWire_46_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_46_T_2 = _ramWire_0_T | _ramWire_46_T_1; // @[mem.scala 25:55]
  wire  _ramWire_46_T_5 = cen & wen & io_memIO_addr == 6'h2e; // @[mem.scala 25:98]
  reg [127:0] ramWire_47_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_47_T_1 = ramWire_47_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_47_T_2 = _ramWire_0_T | _ramWire_47_T_1; // @[mem.scala 25:55]
  wire  _ramWire_47_T_5 = cen & wen & io_memIO_addr == 6'h2f; // @[mem.scala 25:98]
  reg [127:0] ramWire_48_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_48_T_1 = ramWire_48_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_48_T_2 = _ramWire_0_T | _ramWire_48_T_1; // @[mem.scala 25:55]
  wire  _ramWire_48_T_5 = cen & wen & io_memIO_addr == 6'h30; // @[mem.scala 25:98]
  reg [127:0] ramWire_49_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_49_T_1 = ramWire_49_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_49_T_2 = _ramWire_0_T | _ramWire_49_T_1; // @[mem.scala 25:55]
  wire  _ramWire_49_T_5 = cen & wen & io_memIO_addr == 6'h31; // @[mem.scala 25:98]
  reg [127:0] ramWire_50_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_50_T_1 = ramWire_50_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_50_T_2 = _ramWire_0_T | _ramWire_50_T_1; // @[mem.scala 25:55]
  wire  _ramWire_50_T_5 = cen & wen & io_memIO_addr == 6'h32; // @[mem.scala 25:98]
  reg [127:0] ramWire_51_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_51_T_1 = ramWire_51_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_51_T_2 = _ramWire_0_T | _ramWire_51_T_1; // @[mem.scala 25:55]
  wire  _ramWire_51_T_5 = cen & wen & io_memIO_addr == 6'h33; // @[mem.scala 25:98]
  reg [127:0] ramWire_52_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_52_T_1 = ramWire_52_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_52_T_2 = _ramWire_0_T | _ramWire_52_T_1; // @[mem.scala 25:55]
  wire  _ramWire_52_T_5 = cen & wen & io_memIO_addr == 6'h34; // @[mem.scala 25:98]
  reg [127:0] ramWire_53_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_53_T_1 = ramWire_53_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_53_T_2 = _ramWire_0_T | _ramWire_53_T_1; // @[mem.scala 25:55]
  wire  _ramWire_53_T_5 = cen & wen & io_memIO_addr == 6'h35; // @[mem.scala 25:98]
  reg [127:0] ramWire_54_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_54_T_1 = ramWire_54_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_54_T_2 = _ramWire_0_T | _ramWire_54_T_1; // @[mem.scala 25:55]
  wire  _ramWire_54_T_5 = cen & wen & io_memIO_addr == 6'h36; // @[mem.scala 25:98]
  reg [127:0] ramWire_55_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_55_T_1 = ramWire_55_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_55_T_2 = _ramWire_0_T | _ramWire_55_T_1; // @[mem.scala 25:55]
  wire  _ramWire_55_T_5 = cen & wen & io_memIO_addr == 6'h37; // @[mem.scala 25:98]
  reg [127:0] ramWire_56_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_56_T_1 = ramWire_56_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_56_T_2 = _ramWire_0_T | _ramWire_56_T_1; // @[mem.scala 25:55]
  wire  _ramWire_56_T_5 = cen & wen & io_memIO_addr == 6'h38; // @[mem.scala 25:98]
  reg [127:0] ramWire_57_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_57_T_1 = ramWire_57_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_57_T_2 = _ramWire_0_T | _ramWire_57_T_1; // @[mem.scala 25:55]
  wire  _ramWire_57_T_5 = cen & wen & io_memIO_addr == 6'h39; // @[mem.scala 25:98]
  reg [127:0] ramWire_58_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_58_T_1 = ramWire_58_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_58_T_2 = _ramWire_0_T | _ramWire_58_T_1; // @[mem.scala 25:55]
  wire  _ramWire_58_T_5 = cen & wen & io_memIO_addr == 6'h3a; // @[mem.scala 25:98]
  reg [127:0] ramWire_59_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_59_T_1 = ramWire_59_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_59_T_2 = _ramWire_0_T | _ramWire_59_T_1; // @[mem.scala 25:55]
  wire  _ramWire_59_T_5 = cen & wen & io_memIO_addr == 6'h3b; // @[mem.scala 25:98]
  reg [127:0] ramWire_60_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_60_T_1 = ramWire_60_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_60_T_2 = _ramWire_0_T | _ramWire_60_T_1; // @[mem.scala 25:55]
  wire  _ramWire_60_T_5 = cen & wen & io_memIO_addr == 6'h3c; // @[mem.scala 25:98]
  reg [127:0] ramWire_61_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_61_T_1 = ramWire_61_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_61_T_2 = _ramWire_0_T | _ramWire_61_T_1; // @[mem.scala 25:55]
  wire  _ramWire_61_T_5 = cen & wen & io_memIO_addr == 6'h3d; // @[mem.scala 25:98]
  reg [127:0] ramWire_62_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_62_T_1 = ramWire_62_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_62_T_2 = _ramWire_0_T | _ramWire_62_T_1; // @[mem.scala 25:55]
  wire  _ramWire_62_T_5 = cen & wen & io_memIO_addr == 6'h3e; // @[mem.scala 25:98]
  reg [127:0] ramWire_63_r; // @[Reg.scala 15:16]
  wire [127:0] _ramWire_63_T_1 = ramWire_63_r & io_memIO_wmask; // @[mem.scala 25:69]
  wire [127:0] _ramWire_63_T_2 = _ramWire_0_T | _ramWire_63_T_1; // @[mem.scala 25:55]
  wire  _ramWire_63_T_5 = cen & wen & io_memIO_addr == 6'h3f; // @[mem.scala 25:98]
  wire [127:0] _io_memIO_rdata_T_1 = 6'h1 == io_memIO_addr ? ramWire_1_r : ramWire_0_r; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_3 = 6'h2 == io_memIO_addr ? ramWire_2_r : _io_memIO_rdata_T_1; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_5 = 6'h3 == io_memIO_addr ? ramWire_3_r : _io_memIO_rdata_T_3; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_7 = 6'h4 == io_memIO_addr ? ramWire_4_r : _io_memIO_rdata_T_5; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_9 = 6'h5 == io_memIO_addr ? ramWire_5_r : _io_memIO_rdata_T_7; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_11 = 6'h6 == io_memIO_addr ? ramWire_6_r : _io_memIO_rdata_T_9; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_13 = 6'h7 == io_memIO_addr ? ramWire_7_r : _io_memIO_rdata_T_11; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_15 = 6'h8 == io_memIO_addr ? ramWire_8_r : _io_memIO_rdata_T_13; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_17 = 6'h9 == io_memIO_addr ? ramWire_9_r : _io_memIO_rdata_T_15; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_19 = 6'ha == io_memIO_addr ? ramWire_10_r : _io_memIO_rdata_T_17; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_21 = 6'hb == io_memIO_addr ? ramWire_11_r : _io_memIO_rdata_T_19; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_23 = 6'hc == io_memIO_addr ? ramWire_12_r : _io_memIO_rdata_T_21; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_25 = 6'hd == io_memIO_addr ? ramWire_13_r : _io_memIO_rdata_T_23; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_27 = 6'he == io_memIO_addr ? ramWire_14_r : _io_memIO_rdata_T_25; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_29 = 6'hf == io_memIO_addr ? ramWire_15_r : _io_memIO_rdata_T_27; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_31 = 6'h10 == io_memIO_addr ? ramWire_16_r : _io_memIO_rdata_T_29; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_33 = 6'h11 == io_memIO_addr ? ramWire_17_r : _io_memIO_rdata_T_31; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_35 = 6'h12 == io_memIO_addr ? ramWire_18_r : _io_memIO_rdata_T_33; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_37 = 6'h13 == io_memIO_addr ? ramWire_19_r : _io_memIO_rdata_T_35; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_39 = 6'h14 == io_memIO_addr ? ramWire_20_r : _io_memIO_rdata_T_37; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_41 = 6'h15 == io_memIO_addr ? ramWire_21_r : _io_memIO_rdata_T_39; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_43 = 6'h16 == io_memIO_addr ? ramWire_22_r : _io_memIO_rdata_T_41; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_45 = 6'h17 == io_memIO_addr ? ramWire_23_r : _io_memIO_rdata_T_43; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_47 = 6'h18 == io_memIO_addr ? ramWire_24_r : _io_memIO_rdata_T_45; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_49 = 6'h19 == io_memIO_addr ? ramWire_25_r : _io_memIO_rdata_T_47; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_51 = 6'h1a == io_memIO_addr ? ramWire_26_r : _io_memIO_rdata_T_49; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_53 = 6'h1b == io_memIO_addr ? ramWire_27_r : _io_memIO_rdata_T_51; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_55 = 6'h1c == io_memIO_addr ? ramWire_28_r : _io_memIO_rdata_T_53; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_57 = 6'h1d == io_memIO_addr ? ramWire_29_r : _io_memIO_rdata_T_55; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_59 = 6'h1e == io_memIO_addr ? ramWire_30_r : _io_memIO_rdata_T_57; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_61 = 6'h1f == io_memIO_addr ? ramWire_31_r : _io_memIO_rdata_T_59; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_63 = 6'h20 == io_memIO_addr ? ramWire_32_r : _io_memIO_rdata_T_61; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_65 = 6'h21 == io_memIO_addr ? ramWire_33_r : _io_memIO_rdata_T_63; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_67 = 6'h22 == io_memIO_addr ? ramWire_34_r : _io_memIO_rdata_T_65; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_69 = 6'h23 == io_memIO_addr ? ramWire_35_r : _io_memIO_rdata_T_67; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_71 = 6'h24 == io_memIO_addr ? ramWire_36_r : _io_memIO_rdata_T_69; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_73 = 6'h25 == io_memIO_addr ? ramWire_37_r : _io_memIO_rdata_T_71; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_75 = 6'h26 == io_memIO_addr ? ramWire_38_r : _io_memIO_rdata_T_73; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_77 = 6'h27 == io_memIO_addr ? ramWire_39_r : _io_memIO_rdata_T_75; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_79 = 6'h28 == io_memIO_addr ? ramWire_40_r : _io_memIO_rdata_T_77; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_81 = 6'h29 == io_memIO_addr ? ramWire_41_r : _io_memIO_rdata_T_79; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_83 = 6'h2a == io_memIO_addr ? ramWire_42_r : _io_memIO_rdata_T_81; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_85 = 6'h2b == io_memIO_addr ? ramWire_43_r : _io_memIO_rdata_T_83; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_87 = 6'h2c == io_memIO_addr ? ramWire_44_r : _io_memIO_rdata_T_85; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_89 = 6'h2d == io_memIO_addr ? ramWire_45_r : _io_memIO_rdata_T_87; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_91 = 6'h2e == io_memIO_addr ? ramWire_46_r : _io_memIO_rdata_T_89; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_93 = 6'h2f == io_memIO_addr ? ramWire_47_r : _io_memIO_rdata_T_91; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_95 = 6'h30 == io_memIO_addr ? ramWire_48_r : _io_memIO_rdata_T_93; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_97 = 6'h31 == io_memIO_addr ? ramWire_49_r : _io_memIO_rdata_T_95; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_99 = 6'h32 == io_memIO_addr ? ramWire_50_r : _io_memIO_rdata_T_97; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_101 = 6'h33 == io_memIO_addr ? ramWire_51_r : _io_memIO_rdata_T_99; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_103 = 6'h34 == io_memIO_addr ? ramWire_52_r : _io_memIO_rdata_T_101; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_105 = 6'h35 == io_memIO_addr ? ramWire_53_r : _io_memIO_rdata_T_103; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_107 = 6'h36 == io_memIO_addr ? ramWire_54_r : _io_memIO_rdata_T_105; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_109 = 6'h37 == io_memIO_addr ? ramWire_55_r : _io_memIO_rdata_T_107; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_111 = 6'h38 == io_memIO_addr ? ramWire_56_r : _io_memIO_rdata_T_109; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_113 = 6'h39 == io_memIO_addr ? ramWire_57_r : _io_memIO_rdata_T_111; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_115 = 6'h3a == io_memIO_addr ? ramWire_58_r : _io_memIO_rdata_T_113; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_117 = 6'h3b == io_memIO_addr ? ramWire_59_r : _io_memIO_rdata_T_115; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_119 = 6'h3c == io_memIO_addr ? ramWire_60_r : _io_memIO_rdata_T_117; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_121 = 6'h3d == io_memIO_addr ? ramWire_61_r : _io_memIO_rdata_T_119; // @[Mux.scala 80:57]
  wire [127:0] _io_memIO_rdata_T_123 = 6'h3e == io_memIO_addr ? ramWire_62_r : _io_memIO_rdata_T_121; // @[Mux.scala 80:57]
  assign io_memIO_rdata = 6'h3f == io_memIO_addr ? ramWire_63_r : _io_memIO_rdata_T_123; // @[Mux.scala 80:57]
  always @(posedge clock) begin
    if (_ramWire_0_T_5) begin // @[Reg.scala 16:19]
      ramWire_0_r <= _ramWire_0_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_1_T_5) begin // @[Reg.scala 16:19]
      ramWire_1_r <= _ramWire_1_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_2_T_5) begin // @[Reg.scala 16:19]
      ramWire_2_r <= _ramWire_2_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_3_T_5) begin // @[Reg.scala 16:19]
      ramWire_3_r <= _ramWire_3_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_4_T_5) begin // @[Reg.scala 16:19]
      ramWire_4_r <= _ramWire_4_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_5_T_5) begin // @[Reg.scala 16:19]
      ramWire_5_r <= _ramWire_5_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_6_T_5) begin // @[Reg.scala 16:19]
      ramWire_6_r <= _ramWire_6_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_7_T_5) begin // @[Reg.scala 16:19]
      ramWire_7_r <= _ramWire_7_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_8_T_5) begin // @[Reg.scala 16:19]
      ramWire_8_r <= _ramWire_8_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_9_T_5) begin // @[Reg.scala 16:19]
      ramWire_9_r <= _ramWire_9_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_10_T_5) begin // @[Reg.scala 16:19]
      ramWire_10_r <= _ramWire_10_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_11_T_5) begin // @[Reg.scala 16:19]
      ramWire_11_r <= _ramWire_11_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_12_T_5) begin // @[Reg.scala 16:19]
      ramWire_12_r <= _ramWire_12_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_13_T_5) begin // @[Reg.scala 16:19]
      ramWire_13_r <= _ramWire_13_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_14_T_5) begin // @[Reg.scala 16:19]
      ramWire_14_r <= _ramWire_14_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_15_T_5) begin // @[Reg.scala 16:19]
      ramWire_15_r <= _ramWire_15_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_16_T_5) begin // @[Reg.scala 16:19]
      ramWire_16_r <= _ramWire_16_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_17_T_5) begin // @[Reg.scala 16:19]
      ramWire_17_r <= _ramWire_17_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_18_T_5) begin // @[Reg.scala 16:19]
      ramWire_18_r <= _ramWire_18_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_19_T_5) begin // @[Reg.scala 16:19]
      ramWire_19_r <= _ramWire_19_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_20_T_5) begin // @[Reg.scala 16:19]
      ramWire_20_r <= _ramWire_20_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_21_T_5) begin // @[Reg.scala 16:19]
      ramWire_21_r <= _ramWire_21_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_22_T_5) begin // @[Reg.scala 16:19]
      ramWire_22_r <= _ramWire_22_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_23_T_5) begin // @[Reg.scala 16:19]
      ramWire_23_r <= _ramWire_23_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_24_T_5) begin // @[Reg.scala 16:19]
      ramWire_24_r <= _ramWire_24_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_25_T_5) begin // @[Reg.scala 16:19]
      ramWire_25_r <= _ramWire_25_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_26_T_5) begin // @[Reg.scala 16:19]
      ramWire_26_r <= _ramWire_26_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_27_T_5) begin // @[Reg.scala 16:19]
      ramWire_27_r <= _ramWire_27_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_28_T_5) begin // @[Reg.scala 16:19]
      ramWire_28_r <= _ramWire_28_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_29_T_5) begin // @[Reg.scala 16:19]
      ramWire_29_r <= _ramWire_29_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_30_T_5) begin // @[Reg.scala 16:19]
      ramWire_30_r <= _ramWire_30_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_31_T_5) begin // @[Reg.scala 16:19]
      ramWire_31_r <= _ramWire_31_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_32_T_5) begin // @[Reg.scala 16:19]
      ramWire_32_r <= _ramWire_32_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_33_T_5) begin // @[Reg.scala 16:19]
      ramWire_33_r <= _ramWire_33_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_34_T_5) begin // @[Reg.scala 16:19]
      ramWire_34_r <= _ramWire_34_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_35_T_5) begin // @[Reg.scala 16:19]
      ramWire_35_r <= _ramWire_35_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_36_T_5) begin // @[Reg.scala 16:19]
      ramWire_36_r <= _ramWire_36_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_37_T_5) begin // @[Reg.scala 16:19]
      ramWire_37_r <= _ramWire_37_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_38_T_5) begin // @[Reg.scala 16:19]
      ramWire_38_r <= _ramWire_38_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_39_T_5) begin // @[Reg.scala 16:19]
      ramWire_39_r <= _ramWire_39_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_40_T_5) begin // @[Reg.scala 16:19]
      ramWire_40_r <= _ramWire_40_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_41_T_5) begin // @[Reg.scala 16:19]
      ramWire_41_r <= _ramWire_41_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_42_T_5) begin // @[Reg.scala 16:19]
      ramWire_42_r <= _ramWire_42_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_43_T_5) begin // @[Reg.scala 16:19]
      ramWire_43_r <= _ramWire_43_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_44_T_5) begin // @[Reg.scala 16:19]
      ramWire_44_r <= _ramWire_44_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_45_T_5) begin // @[Reg.scala 16:19]
      ramWire_45_r <= _ramWire_45_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_46_T_5) begin // @[Reg.scala 16:19]
      ramWire_46_r <= _ramWire_46_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_47_T_5) begin // @[Reg.scala 16:19]
      ramWire_47_r <= _ramWire_47_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_48_T_5) begin // @[Reg.scala 16:19]
      ramWire_48_r <= _ramWire_48_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_49_T_5) begin // @[Reg.scala 16:19]
      ramWire_49_r <= _ramWire_49_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_50_T_5) begin // @[Reg.scala 16:19]
      ramWire_50_r <= _ramWire_50_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_51_T_5) begin // @[Reg.scala 16:19]
      ramWire_51_r <= _ramWire_51_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_52_T_5) begin // @[Reg.scala 16:19]
      ramWire_52_r <= _ramWire_52_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_53_T_5) begin // @[Reg.scala 16:19]
      ramWire_53_r <= _ramWire_53_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_54_T_5) begin // @[Reg.scala 16:19]
      ramWire_54_r <= _ramWire_54_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_55_T_5) begin // @[Reg.scala 16:19]
      ramWire_55_r <= _ramWire_55_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_56_T_5) begin // @[Reg.scala 16:19]
      ramWire_56_r <= _ramWire_56_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_57_T_5) begin // @[Reg.scala 16:19]
      ramWire_57_r <= _ramWire_57_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_58_T_5) begin // @[Reg.scala 16:19]
      ramWire_58_r <= _ramWire_58_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_59_T_5) begin // @[Reg.scala 16:19]
      ramWire_59_r <= _ramWire_59_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_60_T_5) begin // @[Reg.scala 16:19]
      ramWire_60_r <= _ramWire_60_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_61_T_5) begin // @[Reg.scala 16:19]
      ramWire_61_r <= _ramWire_61_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_62_T_5) begin // @[Reg.scala 16:19]
      ramWire_62_r <= _ramWire_62_T_2; // @[Reg.scala 16:23]
    end
    if (_ramWire_63_T_5) begin // @[Reg.scala 16:19]
      ramWire_63_r <= _ramWire_63_T_2; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  ramWire_0_r = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  ramWire_1_r = _RAND_1[127:0];
  _RAND_2 = {4{`RANDOM}};
  ramWire_2_r = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  ramWire_3_r = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  ramWire_4_r = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  ramWire_5_r = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  ramWire_6_r = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  ramWire_7_r = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  ramWire_8_r = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  ramWire_9_r = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  ramWire_10_r = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  ramWire_11_r = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  ramWire_12_r = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  ramWire_13_r = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  ramWire_14_r = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  ramWire_15_r = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  ramWire_16_r = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  ramWire_17_r = _RAND_17[127:0];
  _RAND_18 = {4{`RANDOM}};
  ramWire_18_r = _RAND_18[127:0];
  _RAND_19 = {4{`RANDOM}};
  ramWire_19_r = _RAND_19[127:0];
  _RAND_20 = {4{`RANDOM}};
  ramWire_20_r = _RAND_20[127:0];
  _RAND_21 = {4{`RANDOM}};
  ramWire_21_r = _RAND_21[127:0];
  _RAND_22 = {4{`RANDOM}};
  ramWire_22_r = _RAND_22[127:0];
  _RAND_23 = {4{`RANDOM}};
  ramWire_23_r = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  ramWire_24_r = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  ramWire_25_r = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  ramWire_26_r = _RAND_26[127:0];
  _RAND_27 = {4{`RANDOM}};
  ramWire_27_r = _RAND_27[127:0];
  _RAND_28 = {4{`RANDOM}};
  ramWire_28_r = _RAND_28[127:0];
  _RAND_29 = {4{`RANDOM}};
  ramWire_29_r = _RAND_29[127:0];
  _RAND_30 = {4{`RANDOM}};
  ramWire_30_r = _RAND_30[127:0];
  _RAND_31 = {4{`RANDOM}};
  ramWire_31_r = _RAND_31[127:0];
  _RAND_32 = {4{`RANDOM}};
  ramWire_32_r = _RAND_32[127:0];
  _RAND_33 = {4{`RANDOM}};
  ramWire_33_r = _RAND_33[127:0];
  _RAND_34 = {4{`RANDOM}};
  ramWire_34_r = _RAND_34[127:0];
  _RAND_35 = {4{`RANDOM}};
  ramWire_35_r = _RAND_35[127:0];
  _RAND_36 = {4{`RANDOM}};
  ramWire_36_r = _RAND_36[127:0];
  _RAND_37 = {4{`RANDOM}};
  ramWire_37_r = _RAND_37[127:0];
  _RAND_38 = {4{`RANDOM}};
  ramWire_38_r = _RAND_38[127:0];
  _RAND_39 = {4{`RANDOM}};
  ramWire_39_r = _RAND_39[127:0];
  _RAND_40 = {4{`RANDOM}};
  ramWire_40_r = _RAND_40[127:0];
  _RAND_41 = {4{`RANDOM}};
  ramWire_41_r = _RAND_41[127:0];
  _RAND_42 = {4{`RANDOM}};
  ramWire_42_r = _RAND_42[127:0];
  _RAND_43 = {4{`RANDOM}};
  ramWire_43_r = _RAND_43[127:0];
  _RAND_44 = {4{`RANDOM}};
  ramWire_44_r = _RAND_44[127:0];
  _RAND_45 = {4{`RANDOM}};
  ramWire_45_r = _RAND_45[127:0];
  _RAND_46 = {4{`RANDOM}};
  ramWire_46_r = _RAND_46[127:0];
  _RAND_47 = {4{`RANDOM}};
  ramWire_47_r = _RAND_47[127:0];
  _RAND_48 = {4{`RANDOM}};
  ramWire_48_r = _RAND_48[127:0];
  _RAND_49 = {4{`RANDOM}};
  ramWire_49_r = _RAND_49[127:0];
  _RAND_50 = {4{`RANDOM}};
  ramWire_50_r = _RAND_50[127:0];
  _RAND_51 = {4{`RANDOM}};
  ramWire_51_r = _RAND_51[127:0];
  _RAND_52 = {4{`RANDOM}};
  ramWire_52_r = _RAND_52[127:0];
  _RAND_53 = {4{`RANDOM}};
  ramWire_53_r = _RAND_53[127:0];
  _RAND_54 = {4{`RANDOM}};
  ramWire_54_r = _RAND_54[127:0];
  _RAND_55 = {4{`RANDOM}};
  ramWire_55_r = _RAND_55[127:0];
  _RAND_56 = {4{`RANDOM}};
  ramWire_56_r = _RAND_56[127:0];
  _RAND_57 = {4{`RANDOM}};
  ramWire_57_r = _RAND_57[127:0];
  _RAND_58 = {4{`RANDOM}};
  ramWire_58_r = _RAND_58[127:0];
  _RAND_59 = {4{`RANDOM}};
  ramWire_59_r = _RAND_59[127:0];
  _RAND_60 = {4{`RANDOM}};
  ramWire_60_r = _RAND_60[127:0];
  _RAND_61 = {4{`RANDOM}};
  ramWire_61_r = _RAND_61[127:0];
  _RAND_62 = {4{`RANDOM}};
  ramWire_62_r = _RAND_62[127:0];
  _RAND_63 = {4{`RANDOM}};
  ramWire_63_r = _RAND_63[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_041728(
  input         clock,
  input         reset,
  input         io_dmaster_awready,
  output        io_dmaster_awvalid,
  output [3:0]  io_dmaster_awid,
  output [31:0] io_dmaster_awaddr,
  output [7:0]  io_dmaster_awlen,
  output [2:0]  io_dmaster_awsize,
  output [1:0]  io_dmaster_awburst,
  input         io_dmaster_wready,
  output        io_dmaster_wvalid,
  output [63:0] io_dmaster_wdata,
  output [7:0]  io_dmaster_wstrb,
  output        io_dmaster_wlast,
  output        io_dmaster_bready,
  input         io_dmaster_bvalid,
  input  [3:0]  io_dmaster_bid,
  input  [1:0]  io_dmaster_bresp,
  input         io_dmaster_arready,
  output        io_dmaster_arvalid,
  output [3:0]  io_dmaster_arid,
  output [31:0] io_dmaster_araddr,
  output [7:0]  io_dmaster_arlen,
  output [2:0]  io_dmaster_arsize,
  output [1:0]  io_dmaster_arburst,
  output        io_dmaster_rready,
  input         io_dmaster_rvalid,
  input  [3:0]  io_dmaster_rid,
  input  [1:0]  io_dmaster_rresp,
  input  [63:0] io_dmaster_rdata,
  input         io_dmaster_rlast,
  output        io_mmio_valid,
  input         io_mmio_ready,
  input  [63:0] io_mmio_data_read,
  output [63:0] io_mmio_data_write,
  output        io_mmio_wen,
  output [31:0] io_mmio_addr,
  output [1:0]  io_mmio_rsize,
  output [7:0]  io_mmio_mask
);
  wire  dmaIns_clock; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_reset; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataIn_arready; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataIn_arvalid; // @[ysyx_22041728.scala 29:22]
  wire [31:0] dmaIns_io_dataIn_araddr; // @[ysyx_22041728.scala 29:22]
  wire [7:0] dmaIns_io_dataIn_arlen; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataIn_rready; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataIn_rvalid; // @[ysyx_22041728.scala 29:22]
  wire [63:0] dmaIns_io_dataIn_rdata; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataIn_rlast; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataOutMMIO_valid; // @[ysyx_22041728.scala 29:22]
  wire [63:0] dmaIns_io_dataOutMMIO_data_write; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_io_dataOutMMIO_wen; // @[ysyx_22041728.scala 29:22]
  wire [31:0] dmaIns_io_dataOutMMIO_addr; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_dmaEn_0; // @[ysyx_22041728.scala 29:22]
  wire [191:0] dmaIns_dmaCtrl_0; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_blockDMA_0; // @[ysyx_22041728.scala 29:22]
  wire  dmaIns_DMABuzy_0; // @[ysyx_22041728.scala 29:22]
  wire  riscvIns_clock; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_reset; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_io_instIO_valid; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_io_instIO_ready; // @[ysyx_22041728.scala 31:24]
  wire [63:0] riscvIns_io_instIO_data_read; // @[ysyx_22041728.scala 31:24]
  wire [31:0] riscvIns_io_instIO_addr; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_io_dataIO_valid; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_io_dataIO_ready; // @[ysyx_22041728.scala 31:24]
  wire [63:0] riscvIns_io_dataIO_data_read; // @[ysyx_22041728.scala 31:24]
  wire [63:0] riscvIns_io_dataIO_data_write; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_io_dataIO_wen; // @[ysyx_22041728.scala 31:24]
  wire [31:0] riscvIns_io_dataIO_addr; // @[ysyx_22041728.scala 31:24]
  wire [1:0] riscvIns_io_dataIO_rsize; // @[ysyx_22041728.scala 31:24]
  wire [7:0] riscvIns_io_dataIO_mask; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_dmaEn_0; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_intrTimeCnt_0; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_startTimeCnt; // @[ysyx_22041728.scala 31:24]
  wire [191:0] riscvIns_dmaCtrl; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_blockDMA_0; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_block2_0; // @[ysyx_22041728.scala 31:24]
  wire  riscvIns_fencei_0; // @[ysyx_22041728.scala 31:24]
  wire  iCache_clock; // @[ysyx_22041728.scala 32:22]
  wire  iCache_reset; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 32:22]
  wire [31:0] iCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 32:22]
  wire [7:0] iCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_cacheOut_r_valid_i; // @[ysyx_22041728.scala 32:22]
  wire [63:0] iCache_io_cacheOut_r_data_i; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_cacheOut_r_last_i; // @[ysyx_22041728.scala 32:22]
  wire [31:0] iCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_cacheIn_valid; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_cacheIn_ready; // @[ysyx_22041728.scala 32:22]
  wire [63:0] iCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 32:22]
  wire [31:0] iCache_io_cacheIn_addr; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 32:22]
  wire [5:0] iCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_0_rdata; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 32:22]
  wire [5:0] iCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_1_rdata; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 32:22]
  wire [5:0] iCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_2_rdata; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 32:22]
  wire  iCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 32:22]
  wire [5:0] iCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 32:22]
  wire [127:0] iCache_io_SRAMIO_3_rdata; // @[ysyx_22041728.scala 32:22]
  wire  iCache_updataICache_0; // @[ysyx_22041728.scala 32:22]
  wire  axiIIO_clock; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_reset; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_awready; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 34:22]
  wire [31:0] axiIIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 34:22]
  wire [2:0] axiIIO_io_axiIO_awsize; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_wready; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 34:22]
  wire [63:0] axiIIO_io_axiIO_wdata; // @[ysyx_22041728.scala 34:22]
  wire [7:0] axiIIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_wlast; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_bready; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_bvalid; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_arready; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 34:22]
  wire [31:0] axiIIO_io_axiIO_araddr; // @[ysyx_22041728.scala 34:22]
  wire [7:0] axiIIO_io_axiIO_arlen; // @[ysyx_22041728.scala 34:22]
  wire [2:0] axiIIO_io_axiIO_arsize; // @[ysyx_22041728.scala 34:22]
  wire [1:0] axiIIO_io_axiIO_arburst; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_rready; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_rvalid; // @[ysyx_22041728.scala 34:22]
  wire [63:0] axiIIO_io_axiIO_rdata; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_axiIO_rlast; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_cache_ar_valid_o; // @[ysyx_22041728.scala 34:22]
  wire [31:0] axiIIO_io_cache_ar_addr_o; // @[ysyx_22041728.scala 34:22]
  wire [7:0] axiIIO_io_cache_ar_len_o; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 34:22]
  wire [63:0] axiIIO_io_cache_r_data_i; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_cache_r_last_i; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_cache_w_valid_o; // @[ysyx_22041728.scala 34:22]
  wire  axiIIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 34:22]
  wire [63:0] axiIIO_io_cache_w_data_o; // @[ysyx_22041728.scala 34:22]
  wire [31:0] axiIIO_io_cache_w_addr_o; // @[ysyx_22041728.scala 34:22]
  wire [7:0] axiIIO_io_cache_w_mask_o; // @[ysyx_22041728.scala 34:22]
  wire [1:0] axiIIO_io_cache_wsize; // @[ysyx_22041728.scala 34:22]
  wire  dArbIns_io_arbIn_valid; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbIn_ready; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbIn_data_read; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbIn_data_write; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbIn_wen; // @[ysyx_22041728.scala 37:23]
  wire [31:0] dArbIns_io_arbIn_addr; // @[ysyx_22041728.scala 37:23]
  wire [1:0] dArbIns_io_arbIn_rsize; // @[ysyx_22041728.scala 37:23]
  wire [7:0] dArbIns_io_arbIn_mask; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbMMIO_valid; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbMMIO_ready; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbMMIO_data_read; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbMMIO_data_write; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbMMIO_wen; // @[ysyx_22041728.scala 37:23]
  wire [31:0] dArbIns_io_arbMMIO_addr; // @[ysyx_22041728.scala 37:23]
  wire [1:0] dArbIns_io_arbMMIO_rsize; // @[ysyx_22041728.scala 37:23]
  wire [7:0] dArbIns_io_arbMMIO_mask; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbClint_valid; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbClint_data_read; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbClint_data_write; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbClint_wen; // @[ysyx_22041728.scala 37:23]
  wire [31:0] dArbIns_io_arbClint_addr; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbDCache_valid; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbDCache_ready; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbDCache_data_read; // @[ysyx_22041728.scala 37:23]
  wire [63:0] dArbIns_io_arbDCache_data_write; // @[ysyx_22041728.scala 37:23]
  wire  dArbIns_io_arbDCache_wen; // @[ysyx_22041728.scala 37:23]
  wire [31:0] dArbIns_io_arbDCache_addr; // @[ysyx_22041728.scala 37:23]
  wire [1:0] dArbIns_io_arbDCache_rsize; // @[ysyx_22041728.scala 37:23]
  wire [7:0] dArbIns_io_arbDCache_mask; // @[ysyx_22041728.scala 37:23]
  wire  mmioDCache_clock; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_reset; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_block; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioIn_valid; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioIn_ready; // @[ysyx_22041728.scala 38:26]
  wire [63:0] mmioDCache_io_mmioIn_data_read; // @[ysyx_22041728.scala 38:26]
  wire [63:0] mmioDCache_io_mmioIn_data_write; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioIn_wen; // @[ysyx_22041728.scala 38:26]
  wire [31:0] mmioDCache_io_mmioIn_addr; // @[ysyx_22041728.scala 38:26]
  wire [1:0] mmioDCache_io_mmioIn_rsize; // @[ysyx_22041728.scala 38:26]
  wire [7:0] mmioDCache_io_mmioIn_mask; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioOut_valid; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioOut_ready; // @[ysyx_22041728.scala 38:26]
  wire [63:0] mmioDCache_io_mmioOut_data_read; // @[ysyx_22041728.scala 38:26]
  wire [63:0] mmioDCache_io_mmioOut_data_write; // @[ysyx_22041728.scala 38:26]
  wire  mmioDCache_io_mmioOut_wen; // @[ysyx_22041728.scala 38:26]
  wire [31:0] mmioDCache_io_mmioOut_addr; // @[ysyx_22041728.scala 38:26]
  wire [1:0] mmioDCache_io_mmioOut_rsize; // @[ysyx_22041728.scala 38:26]
  wire [7:0] mmioDCache_io_mmioOut_mask; // @[ysyx_22041728.scala 38:26]
  wire  dCache_clock; // @[ysyx_22041728.scala 39:22]
  wire  dCache_reset; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 39:22]
  wire [31:0] dCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 39:22]
  wire [7:0] dCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheOut_r_valid_i; // @[ysyx_22041728.scala 39:22]
  wire [63:0] dCache_io_cacheOut_r_data_i; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheOut_r_last_i; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheOut_w_valid_o; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheOut_w_ready_i; // @[ysyx_22041728.scala 39:22]
  wire [63:0] dCache_io_cacheOut_w_data_o; // @[ysyx_22041728.scala 39:22]
  wire [31:0] dCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 39:22]
  wire [7:0] dCache_io_cacheOut_w_mask_o; // @[ysyx_22041728.scala 39:22]
  wire [1:0] dCache_io_cacheOut_wsize; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheIn_valid; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheIn_ready; // @[ysyx_22041728.scala 39:22]
  wire [63:0] dCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 39:22]
  wire [63:0] dCache_io_cacheIn_data_write; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_cacheIn_wen; // @[ysyx_22041728.scala 39:22]
  wire [31:0] dCache_io_cacheIn_addr; // @[ysyx_22041728.scala 39:22]
  wire [1:0] dCache_io_cacheIn_rsize; // @[ysyx_22041728.scala 39:22]
  wire [7:0] dCache_io_cacheIn_mask; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 39:22]
  wire [5:0] dCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_0_rdata; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 39:22]
  wire [5:0] dCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_1_rdata; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 39:22]
  wire [5:0] dCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_2_rdata; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 39:22]
  wire [5:0] dCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 39:22]
  wire [127:0] dCache_io_SRAMIO_3_rdata; // @[ysyx_22041728.scala 39:22]
  wire  dCache_io_block; // @[ysyx_22041728.scala 39:22]
  wire  clintIns_clock; // @[ysyx_22041728.scala 40:25]
  wire  clintIns_reset; // @[ysyx_22041728.scala 40:25]
  wire  clintIns_io_clintIO_valid; // @[ysyx_22041728.scala 40:25]
  wire [63:0] clintIns_io_clintIO_data_read; // @[ysyx_22041728.scala 40:25]
  wire [63:0] clintIns_io_clintIO_data_write; // @[ysyx_22041728.scala 40:25]
  wire  clintIns_io_clintIO_wen; // @[ysyx_22041728.scala 40:25]
  wire [31:0] clintIns_io_clintIO_addr; // @[ysyx_22041728.scala 40:25]
  wire  clintIns_intrTimeCnt_0; // @[ysyx_22041728.scala 40:25]
  wire  clintIns_startTimeCnt_0; // @[ysyx_22041728.scala 40:25]
  wire  axiDIO_clock; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_reset; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_awready; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 46:22]
  wire [31:0] axiDIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 46:22]
  wire [2:0] axiDIO_io_axiIO_awsize; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_wready; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 46:22]
  wire [63:0] axiDIO_io_axiIO_wdata; // @[ysyx_22041728.scala 46:22]
  wire [7:0] axiDIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_wlast; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_bready; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_bvalid; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_arready; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 46:22]
  wire [31:0] axiDIO_io_axiIO_araddr; // @[ysyx_22041728.scala 46:22]
  wire [7:0] axiDIO_io_axiIO_arlen; // @[ysyx_22041728.scala 46:22]
  wire [2:0] axiDIO_io_axiIO_arsize; // @[ysyx_22041728.scala 46:22]
  wire [1:0] axiDIO_io_axiIO_arburst; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_rready; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_rvalid; // @[ysyx_22041728.scala 46:22]
  wire [63:0] axiDIO_io_axiIO_rdata; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_axiIO_rlast; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_cache_ar_valid_o; // @[ysyx_22041728.scala 46:22]
  wire [31:0] axiDIO_io_cache_ar_addr_o; // @[ysyx_22041728.scala 46:22]
  wire [7:0] axiDIO_io_cache_ar_len_o; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 46:22]
  wire [63:0] axiDIO_io_cache_r_data_i; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_cache_r_last_i; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_cache_w_valid_o; // @[ysyx_22041728.scala 46:22]
  wire  axiDIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 46:22]
  wire [63:0] axiDIO_io_cache_w_data_o; // @[ysyx_22041728.scala 46:22]
  wire [31:0] axiDIO_io_cache_w_addr_o; // @[ysyx_22041728.scala 46:22]
  wire [7:0] axiDIO_io_cache_w_mask_o; // @[ysyx_22041728.scala 46:22]
  wire [1:0] axiDIO_io_cache_wsize; // @[ysyx_22041728.scala 46:22]
  wire  imem_clock; // @[ysyx_22041728.scala 53:24]
  wire  imem_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  imem_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] imem_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  dmem_clock; // @[ysyx_22041728.scala 54:24]
  wire  dmem_io_memIO_cen; // @[ysyx_22041728.scala 54:24]
  wire  dmem_io_memIO_wen; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_io_memIO_wdata; // @[ysyx_22041728.scala 54:24]
  wire [5:0] dmem_io_memIO_addr; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_io_memIO_wmask; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_io_memIO_rdata; // @[ysyx_22041728.scala 54:24]
  wire  imem_1_clock; // @[ysyx_22041728.scala 53:24]
  wire  imem_1_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  imem_1_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_1_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] imem_1_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_1_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_1_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  dmem_1_clock; // @[ysyx_22041728.scala 54:24]
  wire  dmem_1_io_memIO_cen; // @[ysyx_22041728.scala 54:24]
  wire  dmem_1_io_memIO_wen; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_1_io_memIO_wdata; // @[ysyx_22041728.scala 54:24]
  wire [5:0] dmem_1_io_memIO_addr; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_1_io_memIO_wmask; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_1_io_memIO_rdata; // @[ysyx_22041728.scala 54:24]
  wire  imem_2_clock; // @[ysyx_22041728.scala 53:24]
  wire  imem_2_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  imem_2_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_2_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] imem_2_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_2_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_2_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  dmem_2_clock; // @[ysyx_22041728.scala 54:24]
  wire  dmem_2_io_memIO_cen; // @[ysyx_22041728.scala 54:24]
  wire  dmem_2_io_memIO_wen; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_2_io_memIO_wdata; // @[ysyx_22041728.scala 54:24]
  wire [5:0] dmem_2_io_memIO_addr; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_2_io_memIO_wmask; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_2_io_memIO_rdata; // @[ysyx_22041728.scala 54:24]
  wire  imem_3_clock; // @[ysyx_22041728.scala 53:24]
  wire  imem_3_io_memIO_cen; // @[ysyx_22041728.scala 53:24]
  wire  imem_3_io_memIO_wen; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_3_io_memIO_wdata; // @[ysyx_22041728.scala 53:24]
  wire [5:0] imem_3_io_memIO_addr; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_3_io_memIO_wmask; // @[ysyx_22041728.scala 53:24]
  wire [127:0] imem_3_io_memIO_rdata; // @[ysyx_22041728.scala 53:24]
  wire  dmem_3_clock; // @[ysyx_22041728.scala 54:24]
  wire  dmem_3_io_memIO_cen; // @[ysyx_22041728.scala 54:24]
  wire  dmem_3_io_memIO_wen; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_3_io_memIO_wdata; // @[ysyx_22041728.scala 54:24]
  wire [5:0] dmem_3_io_memIO_addr; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_3_io_memIO_wmask; // @[ysyx_22041728.scala 54:24]
  wire [127:0] dmem_3_io_memIO_rdata; // @[ysyx_22041728.scala 54:24]
  wire  _io_dmaster_awvalid_T_1 = riscvIns_io_instIO_valid & ~riscvIns_io_instIO_ready; // @[ysyx_22041728.scala 249:34]
  wire  _io_dmaster_awvalid_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_awvalid : axiDIO_io_axiIO_awvalid; // @[ysyx_22041728.scala 248:10]
  wire  DMABuzy_0 = dmaIns_DMABuzy_0;
  wire  _io_dmaster_wvalid_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_wvalid : axiDIO_io_axiIO_wvalid; // @[ysyx_22041728.scala 248:10]
  wire  _io_dmaster_wlast_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_wlast : axiDIO_io_axiIO_wlast; // @[ysyx_22041728.scala 248:10]
  wire  _io_dmaster_bready_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_bready : axiDIO_io_axiIO_bready; // @[ysyx_22041728.scala 248:10]
  wire  _io_dmaster_arvalid_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_arvalid : axiDIO_io_axiIO_arvalid; // @[ysyx_22041728.scala 248:10]
  wire  _io_dmaster_rready_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_rready : axiDIO_io_axiIO_rready; // @[ysyx_22041728.scala 248:10]
  wire [2:0] _io_dmaster_awsize_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_awsize : axiDIO_io_axiIO_awsize; // @[ysyx_22041728.scala 248:10]
  wire [31:0] _io_dmaster_awaddr_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_awaddr : axiDIO_io_axiIO_awaddr; // @[ysyx_22041728.scala 248:10]
  wire [31:0] _io_dmaster_araddr_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_araddr : axiDIO_io_axiIO_araddr; // @[ysyx_22041728.scala 248:10]
  wire [63:0] _io_dmaster_wdata_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_wdata : axiDIO_io_axiIO_wdata; // @[ysyx_22041728.scala 248:10]
  wire [7:0] _io_dmaster_wstrb_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_wstrb : axiDIO_io_axiIO_wstrb; // @[ysyx_22041728.scala 248:10]
  wire [7:0] _io_dmaster_arlen_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_arlen : axiDIO_io_axiIO_arlen; // @[ysyx_22041728.scala 248:10]
  wire [2:0] _io_dmaster_arsize_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_arsize : axiDIO_io_axiIO_arsize; // @[ysyx_22041728.scala 248:10]
  wire [1:0] _io_dmaster_arburst_T_2 = _io_dmaster_awvalid_T_1 ? axiIIO_io_axiIO_arburst : axiDIO_io_axiIO_arburst; // @[ysyx_22041728.scala 248:10]
  DMACtrl dmaIns ( // @[ysyx_22041728.scala 29:22]
    .clock(dmaIns_clock),
    .reset(dmaIns_reset),
    .io_dataIn_arready(dmaIns_io_dataIn_arready),
    .io_dataIn_arvalid(dmaIns_io_dataIn_arvalid),
    .io_dataIn_araddr(dmaIns_io_dataIn_araddr),
    .io_dataIn_arlen(dmaIns_io_dataIn_arlen),
    .io_dataIn_rready(dmaIns_io_dataIn_rready),
    .io_dataIn_rvalid(dmaIns_io_dataIn_rvalid),
    .io_dataIn_rdata(dmaIns_io_dataIn_rdata),
    .io_dataIn_rlast(dmaIns_io_dataIn_rlast),
    .io_dataOutMMIO_valid(dmaIns_io_dataOutMMIO_valid),
    .io_dataOutMMIO_data_write(dmaIns_io_dataOutMMIO_data_write),
    .io_dataOutMMIO_wen(dmaIns_io_dataOutMMIO_wen),
    .io_dataOutMMIO_addr(dmaIns_io_dataOutMMIO_addr),
    .dmaEn_0(dmaIns_dmaEn_0),
    .dmaCtrl_0(dmaIns_dmaCtrl_0),
    .blockDMA_0(dmaIns_blockDMA_0),
    .DMABuzy_0(dmaIns_DMABuzy_0)
  );
  riscv riscvIns ( // @[ysyx_22041728.scala 31:24]
    .clock(riscvIns_clock),
    .reset(riscvIns_reset),
    .io_instIO_valid(riscvIns_io_instIO_valid),
    .io_instIO_ready(riscvIns_io_instIO_ready),
    .io_instIO_data_read(riscvIns_io_instIO_data_read),
    .io_instIO_addr(riscvIns_io_instIO_addr),
    .io_dataIO_valid(riscvIns_io_dataIO_valid),
    .io_dataIO_ready(riscvIns_io_dataIO_ready),
    .io_dataIO_data_read(riscvIns_io_dataIO_data_read),
    .io_dataIO_data_write(riscvIns_io_dataIO_data_write),
    .io_dataIO_wen(riscvIns_io_dataIO_wen),
    .io_dataIO_addr(riscvIns_io_dataIO_addr),
    .io_dataIO_rsize(riscvIns_io_dataIO_rsize),
    .io_dataIO_mask(riscvIns_io_dataIO_mask),
    .dmaEn_0(riscvIns_dmaEn_0),
    .intrTimeCnt_0(riscvIns_intrTimeCnt_0),
    .startTimeCnt(riscvIns_startTimeCnt),
    .dmaCtrl(riscvIns_dmaCtrl),
    .blockDMA_0(riscvIns_blockDMA_0),
    .block2_0(riscvIns_block2_0),
    .fencei_0(riscvIns_fencei_0)
  );
  Icache iCache ( // @[ysyx_22041728.scala 32:22]
    .clock(iCache_clock),
    .reset(iCache_reset),
    .io_cacheOut_ar_valid_o(iCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(iCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(iCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(iCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(iCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(iCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_addr_o(iCache_io_cacheOut_w_addr_o),
    .io_cacheIn_valid(iCache_io_cacheIn_valid),
    .io_cacheIn_ready(iCache_io_cacheIn_ready),
    .io_cacheIn_data_read(iCache_io_cacheIn_data_read),
    .io_cacheIn_addr(iCache_io_cacheIn_addr),
    .io_SRAMIO_0_cen(iCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(iCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(iCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(iCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(iCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(iCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(iCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(iCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(iCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(iCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(iCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(iCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(iCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(iCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(iCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(iCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(iCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(iCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(iCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(iCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(iCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(iCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(iCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(iCache_io_SRAMIO_3_rdata),
    .updataICache_0(iCache_updataICache_0)
  );
  AXICache axiIIO ( // @[ysyx_22041728.scala 34:22]
    .clock(axiIIO_clock),
    .reset(axiIIO_reset),
    .io_axiIO_awready(axiIIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiIIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiIIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiIIO_io_axiIO_awsize),
    .io_axiIO_wready(axiIIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiIIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiIIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiIIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiIIO_io_axiIO_wlast),
    .io_axiIO_bready(axiIIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiIIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiIIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiIIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiIIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiIIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiIIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiIIO_io_axiIO_arburst),
    .io_axiIO_rready(axiIIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiIIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiIIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiIIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiIIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiIIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiIIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiIIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiIIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiIIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiIIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiIIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiIIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiIIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiIIO_io_cache_w_mask_o),
    .io_cache_wsize(axiIIO_io_cache_wsize)
  );
  arbCpu2DCache dArbIns ( // @[ysyx_22041728.scala 37:23]
    .io_arbIn_valid(dArbIns_io_arbIn_valid),
    .io_arbIn_ready(dArbIns_io_arbIn_ready),
    .io_arbIn_data_read(dArbIns_io_arbIn_data_read),
    .io_arbIn_data_write(dArbIns_io_arbIn_data_write),
    .io_arbIn_wen(dArbIns_io_arbIn_wen),
    .io_arbIn_addr(dArbIns_io_arbIn_addr),
    .io_arbIn_rsize(dArbIns_io_arbIn_rsize),
    .io_arbIn_mask(dArbIns_io_arbIn_mask),
    .io_arbMMIO_valid(dArbIns_io_arbMMIO_valid),
    .io_arbMMIO_ready(dArbIns_io_arbMMIO_ready),
    .io_arbMMIO_data_read(dArbIns_io_arbMMIO_data_read),
    .io_arbMMIO_data_write(dArbIns_io_arbMMIO_data_write),
    .io_arbMMIO_wen(dArbIns_io_arbMMIO_wen),
    .io_arbMMIO_addr(dArbIns_io_arbMMIO_addr),
    .io_arbMMIO_rsize(dArbIns_io_arbMMIO_rsize),
    .io_arbMMIO_mask(dArbIns_io_arbMMIO_mask),
    .io_arbClint_valid(dArbIns_io_arbClint_valid),
    .io_arbClint_data_read(dArbIns_io_arbClint_data_read),
    .io_arbClint_data_write(dArbIns_io_arbClint_data_write),
    .io_arbClint_wen(dArbIns_io_arbClint_wen),
    .io_arbClint_addr(dArbIns_io_arbClint_addr),
    .io_arbDCache_valid(dArbIns_io_arbDCache_valid),
    .io_arbDCache_ready(dArbIns_io_arbDCache_ready),
    .io_arbDCache_data_read(dArbIns_io_arbDCache_data_read),
    .io_arbDCache_data_write(dArbIns_io_arbDCache_data_write),
    .io_arbDCache_wen(dArbIns_io_arbDCache_wen),
    .io_arbDCache_addr(dArbIns_io_arbDCache_addr),
    .io_arbDCache_rsize(dArbIns_io_arbDCache_rsize),
    .io_arbDCache_mask(dArbIns_io_arbDCache_mask)
  );
  mmioCache mmioDCache ( // @[ysyx_22041728.scala 38:26]
    .clock(mmioDCache_clock),
    .reset(mmioDCache_reset),
    .io_block(mmioDCache_io_block),
    .io_mmioIn_valid(mmioDCache_io_mmioIn_valid),
    .io_mmioIn_ready(mmioDCache_io_mmioIn_ready),
    .io_mmioIn_data_read(mmioDCache_io_mmioIn_data_read),
    .io_mmioIn_data_write(mmioDCache_io_mmioIn_data_write),
    .io_mmioIn_wen(mmioDCache_io_mmioIn_wen),
    .io_mmioIn_addr(mmioDCache_io_mmioIn_addr),
    .io_mmioIn_rsize(mmioDCache_io_mmioIn_rsize),
    .io_mmioIn_mask(mmioDCache_io_mmioIn_mask),
    .io_mmioOut_valid(mmioDCache_io_mmioOut_valid),
    .io_mmioOut_ready(mmioDCache_io_mmioOut_ready),
    .io_mmioOut_data_read(mmioDCache_io_mmioOut_data_read),
    .io_mmioOut_data_write(mmioDCache_io_mmioOut_data_write),
    .io_mmioOut_wen(mmioDCache_io_mmioOut_wen),
    .io_mmioOut_addr(mmioDCache_io_mmioOut_addr),
    .io_mmioOut_rsize(mmioDCache_io_mmioOut_rsize),
    .io_mmioOut_mask(mmioDCache_io_mmioOut_mask)
  );
  Dcache dCache ( // @[ysyx_22041728.scala 39:22]
    .clock(dCache_clock),
    .reset(dCache_reset),
    .io_cacheOut_ar_valid_o(dCache_io_cacheOut_ar_valid_o),
    .io_cacheOut_ar_addr_o(dCache_io_cacheOut_ar_addr_o),
    .io_cacheOut_ar_len_o(dCache_io_cacheOut_ar_len_o),
    .io_cacheOut_r_valid_i(dCache_io_cacheOut_r_valid_i),
    .io_cacheOut_r_data_i(dCache_io_cacheOut_r_data_i),
    .io_cacheOut_r_last_i(dCache_io_cacheOut_r_last_i),
    .io_cacheOut_w_valid_o(dCache_io_cacheOut_w_valid_o),
    .io_cacheOut_w_ready_i(dCache_io_cacheOut_w_ready_i),
    .io_cacheOut_w_data_o(dCache_io_cacheOut_w_data_o),
    .io_cacheOut_w_addr_o(dCache_io_cacheOut_w_addr_o),
    .io_cacheOut_w_mask_o(dCache_io_cacheOut_w_mask_o),
    .io_cacheOut_wsize(dCache_io_cacheOut_wsize),
    .io_cacheIn_valid(dCache_io_cacheIn_valid),
    .io_cacheIn_ready(dCache_io_cacheIn_ready),
    .io_cacheIn_data_read(dCache_io_cacheIn_data_read),
    .io_cacheIn_data_write(dCache_io_cacheIn_data_write),
    .io_cacheIn_wen(dCache_io_cacheIn_wen),
    .io_cacheIn_addr(dCache_io_cacheIn_addr),
    .io_cacheIn_rsize(dCache_io_cacheIn_rsize),
    .io_cacheIn_mask(dCache_io_cacheIn_mask),
    .io_SRAMIO_0_cen(dCache_io_SRAMIO_0_cen),
    .io_SRAMIO_0_wen(dCache_io_SRAMIO_0_wen),
    .io_SRAMIO_0_wdata(dCache_io_SRAMIO_0_wdata),
    .io_SRAMIO_0_addr(dCache_io_SRAMIO_0_addr),
    .io_SRAMIO_0_wmask(dCache_io_SRAMIO_0_wmask),
    .io_SRAMIO_0_rdata(dCache_io_SRAMIO_0_rdata),
    .io_SRAMIO_1_cen(dCache_io_SRAMIO_1_cen),
    .io_SRAMIO_1_wen(dCache_io_SRAMIO_1_wen),
    .io_SRAMIO_1_wdata(dCache_io_SRAMIO_1_wdata),
    .io_SRAMIO_1_addr(dCache_io_SRAMIO_1_addr),
    .io_SRAMIO_1_wmask(dCache_io_SRAMIO_1_wmask),
    .io_SRAMIO_1_rdata(dCache_io_SRAMIO_1_rdata),
    .io_SRAMIO_2_cen(dCache_io_SRAMIO_2_cen),
    .io_SRAMIO_2_wen(dCache_io_SRAMIO_2_wen),
    .io_SRAMIO_2_wdata(dCache_io_SRAMIO_2_wdata),
    .io_SRAMIO_2_addr(dCache_io_SRAMIO_2_addr),
    .io_SRAMIO_2_wmask(dCache_io_SRAMIO_2_wmask),
    .io_SRAMIO_2_rdata(dCache_io_SRAMIO_2_rdata),
    .io_SRAMIO_3_cen(dCache_io_SRAMIO_3_cen),
    .io_SRAMIO_3_wen(dCache_io_SRAMIO_3_wen),
    .io_SRAMIO_3_wdata(dCache_io_SRAMIO_3_wdata),
    .io_SRAMIO_3_addr(dCache_io_SRAMIO_3_addr),
    .io_SRAMIO_3_wmask(dCache_io_SRAMIO_3_wmask),
    .io_SRAMIO_3_rdata(dCache_io_SRAMIO_3_rdata),
    .io_block(dCache_io_block)
  );
  clint clintIns ( // @[ysyx_22041728.scala 40:25]
    .clock(clintIns_clock),
    .reset(clintIns_reset),
    .io_clintIO_valid(clintIns_io_clintIO_valid),
    .io_clintIO_data_read(clintIns_io_clintIO_data_read),
    .io_clintIO_data_write(clintIns_io_clintIO_data_write),
    .io_clintIO_wen(clintIns_io_clintIO_wen),
    .io_clintIO_addr(clintIns_io_clintIO_addr),
    .intrTimeCnt_0(clintIns_intrTimeCnt_0),
    .startTimeCnt_0(clintIns_startTimeCnt_0)
  );
  AXICache axiDIO ( // @[ysyx_22041728.scala 46:22]
    .clock(axiDIO_clock),
    .reset(axiDIO_reset),
    .io_axiIO_awready(axiDIO_io_axiIO_awready),
    .io_axiIO_awvalid(axiDIO_io_axiIO_awvalid),
    .io_axiIO_awaddr(axiDIO_io_axiIO_awaddr),
    .io_axiIO_awsize(axiDIO_io_axiIO_awsize),
    .io_axiIO_wready(axiDIO_io_axiIO_wready),
    .io_axiIO_wvalid(axiDIO_io_axiIO_wvalid),
    .io_axiIO_wdata(axiDIO_io_axiIO_wdata),
    .io_axiIO_wstrb(axiDIO_io_axiIO_wstrb),
    .io_axiIO_wlast(axiDIO_io_axiIO_wlast),
    .io_axiIO_bready(axiDIO_io_axiIO_bready),
    .io_axiIO_bvalid(axiDIO_io_axiIO_bvalid),
    .io_axiIO_arready(axiDIO_io_axiIO_arready),
    .io_axiIO_arvalid(axiDIO_io_axiIO_arvalid),
    .io_axiIO_araddr(axiDIO_io_axiIO_araddr),
    .io_axiIO_arlen(axiDIO_io_axiIO_arlen),
    .io_axiIO_arsize(axiDIO_io_axiIO_arsize),
    .io_axiIO_arburst(axiDIO_io_axiIO_arburst),
    .io_axiIO_rready(axiDIO_io_axiIO_rready),
    .io_axiIO_rvalid(axiDIO_io_axiIO_rvalid),
    .io_axiIO_rdata(axiDIO_io_axiIO_rdata),
    .io_axiIO_rlast(axiDIO_io_axiIO_rlast),
    .io_cache_ar_valid_o(axiDIO_io_cache_ar_valid_o),
    .io_cache_ar_addr_o(axiDIO_io_cache_ar_addr_o),
    .io_cache_ar_len_o(axiDIO_io_cache_ar_len_o),
    .io_cache_r_valid_i(axiDIO_io_cache_r_valid_i),
    .io_cache_r_data_i(axiDIO_io_cache_r_data_i),
    .io_cache_r_last_i(axiDIO_io_cache_r_last_i),
    .io_cache_w_valid_o(axiDIO_io_cache_w_valid_o),
    .io_cache_w_ready_i(axiDIO_io_cache_w_ready_i),
    .io_cache_w_data_o(axiDIO_io_cache_w_data_o),
    .io_cache_w_addr_o(axiDIO_io_cache_w_addr_o),
    .io_cache_w_mask_o(axiDIO_io_cache_w_mask_o),
    .io_cache_wsize(axiDIO_io_cache_wsize)
  );
  mem imem ( // @[ysyx_22041728.scala 53:24]
    .clock(imem_clock),
    .io_memIO_cen(imem_io_memIO_cen),
    .io_memIO_wen(imem_io_memIO_wen),
    .io_memIO_wdata(imem_io_memIO_wdata),
    .io_memIO_addr(imem_io_memIO_addr),
    .io_memIO_wmask(imem_io_memIO_wmask),
    .io_memIO_rdata(imem_io_memIO_rdata)
  );
  mem dmem ( // @[ysyx_22041728.scala 54:24]
    .clock(dmem_clock),
    .io_memIO_cen(dmem_io_memIO_cen),
    .io_memIO_wen(dmem_io_memIO_wen),
    .io_memIO_wdata(dmem_io_memIO_wdata),
    .io_memIO_addr(dmem_io_memIO_addr),
    .io_memIO_wmask(dmem_io_memIO_wmask),
    .io_memIO_rdata(dmem_io_memIO_rdata)
  );
  mem imem_1 ( // @[ysyx_22041728.scala 53:24]
    .clock(imem_1_clock),
    .io_memIO_cen(imem_1_io_memIO_cen),
    .io_memIO_wen(imem_1_io_memIO_wen),
    .io_memIO_wdata(imem_1_io_memIO_wdata),
    .io_memIO_addr(imem_1_io_memIO_addr),
    .io_memIO_wmask(imem_1_io_memIO_wmask),
    .io_memIO_rdata(imem_1_io_memIO_rdata)
  );
  mem dmem_1 ( // @[ysyx_22041728.scala 54:24]
    .clock(dmem_1_clock),
    .io_memIO_cen(dmem_1_io_memIO_cen),
    .io_memIO_wen(dmem_1_io_memIO_wen),
    .io_memIO_wdata(dmem_1_io_memIO_wdata),
    .io_memIO_addr(dmem_1_io_memIO_addr),
    .io_memIO_wmask(dmem_1_io_memIO_wmask),
    .io_memIO_rdata(dmem_1_io_memIO_rdata)
  );
  mem imem_2 ( // @[ysyx_22041728.scala 53:24]
    .clock(imem_2_clock),
    .io_memIO_cen(imem_2_io_memIO_cen),
    .io_memIO_wen(imem_2_io_memIO_wen),
    .io_memIO_wdata(imem_2_io_memIO_wdata),
    .io_memIO_addr(imem_2_io_memIO_addr),
    .io_memIO_wmask(imem_2_io_memIO_wmask),
    .io_memIO_rdata(imem_2_io_memIO_rdata)
  );
  mem dmem_2 ( // @[ysyx_22041728.scala 54:24]
    .clock(dmem_2_clock),
    .io_memIO_cen(dmem_2_io_memIO_cen),
    .io_memIO_wen(dmem_2_io_memIO_wen),
    .io_memIO_wdata(dmem_2_io_memIO_wdata),
    .io_memIO_addr(dmem_2_io_memIO_addr),
    .io_memIO_wmask(dmem_2_io_memIO_wmask),
    .io_memIO_rdata(dmem_2_io_memIO_rdata)
  );
  mem imem_3 ( // @[ysyx_22041728.scala 53:24]
    .clock(imem_3_clock),
    .io_memIO_cen(imem_3_io_memIO_cen),
    .io_memIO_wen(imem_3_io_memIO_wen),
    .io_memIO_wdata(imem_3_io_memIO_wdata),
    .io_memIO_addr(imem_3_io_memIO_addr),
    .io_memIO_wmask(imem_3_io_memIO_wmask),
    .io_memIO_rdata(imem_3_io_memIO_rdata)
  );
  mem dmem_3 ( // @[ysyx_22041728.scala 54:24]
    .clock(dmem_3_clock),
    .io_memIO_cen(dmem_3_io_memIO_cen),
    .io_memIO_wen(dmem_3_io_memIO_wen),
    .io_memIO_wdata(dmem_3_io_memIO_wdata),
    .io_memIO_addr(dmem_3_io_memIO_addr),
    .io_memIO_wmask(dmem_3_io_memIO_wmask),
    .io_memIO_rdata(dmem_3_io_memIO_rdata)
  );
  assign io_dmaster_awvalid = DMABuzy_0 ? 1'h0 : _io_dmaster_awvalid_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_awid = 4'h0; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_awaddr = DMABuzy_0 ? 32'h0 : _io_dmaster_awaddr_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_awlen = 8'h0; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_awsize = DMABuzy_0 ? 3'h0 : _io_dmaster_awsize_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_awburst = DMABuzy_0 ? 2'h0 : 2'h1; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_wvalid = DMABuzy_0 ? 1'h0 : _io_dmaster_wvalid_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_wdata = DMABuzy_0 ? 64'h0 : _io_dmaster_wdata_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_wstrb = DMABuzy_0 ? 8'h0 : _io_dmaster_wstrb_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_wlast = DMABuzy_0 ? 1'h0 : _io_dmaster_wlast_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_bready = DMABuzy_0 ? 1'h0 : _io_dmaster_bready_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_arvalid = DMABuzy_0 ? dmaIns_io_dataIn_arvalid : _io_dmaster_arvalid_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_arid = 4'h0; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_araddr = DMABuzy_0 ? dmaIns_io_dataIn_araddr : _io_dmaster_araddr_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_arlen = DMABuzy_0 ? dmaIns_io_dataIn_arlen : _io_dmaster_arlen_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_arsize = DMABuzy_0 ? 3'h3 : _io_dmaster_arsize_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_arburst = DMABuzy_0 ? 2'h1 : _io_dmaster_arburst_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_dmaster_rready = DMABuzy_0 ? dmaIns_io_dataIn_rready : _io_dmaster_rready_T_2; // @[ysyx_22041728.scala 245:29]
  assign io_mmio_valid = DMABuzy_0 ? dmaIns_io_dataOutMMIO_valid : mmioDCache_io_mmioOut_valid; // @[ysyx_22041728.scala 302:28]
  assign io_mmio_data_write = DMABuzy_0 ? dmaIns_io_dataOutMMIO_data_write : mmioDCache_io_mmioOut_data_write; // @[ysyx_22041728.scala 302:28]
  assign io_mmio_wen = DMABuzy_0 ? dmaIns_io_dataOutMMIO_wen : mmioDCache_io_mmioOut_wen; // @[ysyx_22041728.scala 302:28]
  assign io_mmio_addr = DMABuzy_0 ? dmaIns_io_dataOutMMIO_addr : mmioDCache_io_mmioOut_addr; // @[ysyx_22041728.scala 302:28]
  assign io_mmio_rsize = DMABuzy_0 ? 2'h3 : mmioDCache_io_mmioOut_rsize; // @[ysyx_22041728.scala 302:28]
  assign io_mmio_mask = DMABuzy_0 ? 8'hff : mmioDCache_io_mmioOut_mask; // @[ysyx_22041728.scala 302:28]
  assign dmaIns_clock = clock;
  assign dmaIns_reset = reset;
  assign dmaIns_io_dataIn_arready = io_dmaster_arready; // @[ysyx_22041728.scala 255:21]
  assign dmaIns_io_dataIn_rvalid = io_dmaster_rvalid; // @[ysyx_22041728.scala 255:21]
  assign dmaIns_io_dataIn_rdata = io_dmaster_rdata; // @[ysyx_22041728.scala 255:21]
  assign dmaIns_io_dataIn_rlast = io_dmaster_rlast; // @[ysyx_22041728.scala 255:21]
  assign dmaIns_dmaEn_0 = riscvIns_dmaEn_0;
  assign dmaIns_dmaCtrl_0 = riscvIns_dmaCtrl;
  assign riscvIns_clock = clock;
  assign riscvIns_reset = reset;
  assign riscvIns_io_instIO_ready = iCache_io_cacheIn_ready; // @[ysyx_22041728.scala 33:22]
  assign riscvIns_io_instIO_data_read = iCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 33:22]
  assign riscvIns_io_dataIO_ready = dArbIns_io_arbIn_ready; // @[ysyx_22041728.scala 41:21]
  assign riscvIns_io_dataIO_data_read = dArbIns_io_arbIn_data_read; // @[ysyx_22041728.scala 41:21]
  assign riscvIns_intrTimeCnt_0 = clintIns_intrTimeCnt_0;
  assign riscvIns_blockDMA_0 = dmaIns_blockDMA_0;
  assign iCache_clock = clock;
  assign iCache_reset = reset;
  assign iCache_io_cacheOut_r_valid_i = axiIIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 35:19]
  assign iCache_io_cacheOut_r_data_i = axiIIO_io_cache_r_data_i; // @[ysyx_22041728.scala 35:19]
  assign iCache_io_cacheOut_r_last_i = axiIIO_io_cache_r_last_i; // @[ysyx_22041728.scala 35:19]
  assign iCache_io_cacheIn_valid = riscvIns_io_instIO_valid; // @[ysyx_22041728.scala 33:22]
  assign iCache_io_cacheIn_addr = riscvIns_io_instIO_addr; // @[ysyx_22041728.scala 33:22]
  assign iCache_io_SRAMIO_0_rdata = imem_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign iCache_io_SRAMIO_1_rdata = imem_1_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign iCache_io_SRAMIO_2_rdata = imem_2_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign iCache_io_SRAMIO_3_rdata = imem_3_io_memIO_rdata; // @[ysyx_22041728.scala 55:20]
  assign iCache_updataICache_0 = riscvIns_fencei_0;
  assign axiIIO_clock = clock;
  assign axiIIO_reset = reset;
  assign axiIIO_io_axiIO_awready = io_dmaster_awready; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_wready = io_dmaster_wready; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_bvalid = io_dmaster_bvalid; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_arready = io_dmaster_arready; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_rvalid = io_dmaster_rvalid; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_rdata = io_dmaster_rdata; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_axiIO_rlast = io_dmaster_rlast; // @[ysyx_22041728.scala 257:24]
  assign axiIIO_io_cache_ar_valid_o = iCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_ar_addr_o = iCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_ar_len_o = iCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_w_valid_o = 1'h0; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_w_data_o = 64'h0; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_w_addr_o = iCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_w_mask_o = 8'h0; // @[ysyx_22041728.scala 35:19]
  assign axiIIO_io_cache_wsize = 2'h2; // @[ysyx_22041728.scala 35:19]
  assign dArbIns_io_arbIn_valid = riscvIns_io_dataIO_valid; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbIn_data_write = riscvIns_io_dataIO_data_write; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbIn_wen = riscvIns_io_dataIO_wen; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbIn_addr = riscvIns_io_dataIO_addr; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbIn_rsize = riscvIns_io_dataIO_rsize; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbIn_mask = riscvIns_io_dataIO_mask; // @[ysyx_22041728.scala 41:21]
  assign dArbIns_io_arbMMIO_ready = mmioDCache_io_mmioIn_ready; // @[ysyx_22041728.scala 42:21]
  assign dArbIns_io_arbMMIO_data_read = mmioDCache_io_mmioIn_data_read; // @[ysyx_22041728.scala 42:21]
  assign dArbIns_io_arbClint_data_read = clintIns_io_clintIO_data_read; // @[ysyx_22041728.scala 44:22]
  assign dArbIns_io_arbDCache_ready = dCache_io_cacheIn_ready; // @[ysyx_22041728.scala 43:24]
  assign dArbIns_io_arbDCache_data_read = dCache_io_cacheIn_data_read; // @[ysyx_22041728.scala 43:24]
  assign mmioDCache_clock = clock;
  assign mmioDCache_reset = reset;
  assign mmioDCache_io_block = riscvIns_block2_0; // @[ysyx_22041728.scala 78:20]
  assign mmioDCache_io_mmioIn_valid = dArbIns_io_arbMMIO_valid; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioIn_data_write = dArbIns_io_arbMMIO_data_write; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioIn_wen = dArbIns_io_arbMMIO_wen; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioIn_addr = dArbIns_io_arbMMIO_addr; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioIn_rsize = dArbIns_io_arbMMIO_rsize; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioIn_mask = dArbIns_io_arbMMIO_mask; // @[ysyx_22041728.scala 42:21]
  assign mmioDCache_io_mmioOut_ready = io_mmio_ready; // @[ysyx_22041728.scala 310:25]
  assign mmioDCache_io_mmioOut_data_read = io_mmio_data_read; // @[ysyx_22041728.scala 310:25]
  assign dCache_clock = clock;
  assign dCache_reset = reset;
  assign dCache_io_cacheOut_r_valid_i = axiDIO_io_cache_r_valid_i; // @[ysyx_22041728.scala 48:18]
  assign dCache_io_cacheOut_r_data_i = axiDIO_io_cache_r_data_i; // @[ysyx_22041728.scala 48:18]
  assign dCache_io_cacheOut_r_last_i = axiDIO_io_cache_r_last_i; // @[ysyx_22041728.scala 48:18]
  assign dCache_io_cacheOut_w_ready_i = axiDIO_io_cache_w_ready_i; // @[ysyx_22041728.scala 48:18]
  assign dCache_io_cacheIn_valid = dArbIns_io_arbDCache_valid; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_cacheIn_data_write = dArbIns_io_arbDCache_data_write; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_cacheIn_wen = dArbIns_io_arbDCache_wen; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_cacheIn_addr = dArbIns_io_arbDCache_addr; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_cacheIn_rsize = dArbIns_io_arbDCache_rsize; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_cacheIn_mask = dArbIns_io_arbDCache_mask; // @[ysyx_22041728.scala 43:24]
  assign dCache_io_SRAMIO_0_rdata = dmem_io_memIO_rdata; // @[ysyx_22041728.scala 56:20]
  assign dCache_io_SRAMIO_1_rdata = dmem_1_io_memIO_rdata; // @[ysyx_22041728.scala 56:20]
  assign dCache_io_SRAMIO_2_rdata = dmem_2_io_memIO_rdata; // @[ysyx_22041728.scala 56:20]
  assign dCache_io_SRAMIO_3_rdata = dmem_3_io_memIO_rdata; // @[ysyx_22041728.scala 56:20]
  assign dCache_io_block = riscvIns_block2_0; // @[ysyx_22041728.scala 78:20]
  assign clintIns_clock = clock;
  assign clintIns_reset = reset;
  assign clintIns_io_clintIO_valid = dArbIns_io_arbClint_valid; // @[ysyx_22041728.scala 44:22]
  assign clintIns_io_clintIO_data_write = dArbIns_io_arbClint_data_write; // @[ysyx_22041728.scala 44:22]
  assign clintIns_io_clintIO_wen = dArbIns_io_arbClint_wen; // @[ysyx_22041728.scala 44:22]
  assign clintIns_io_clintIO_addr = dArbIns_io_arbClint_addr; // @[ysyx_22041728.scala 44:22]
  assign clintIns_startTimeCnt_0 = riscvIns_startTimeCnt;
  assign axiDIO_clock = clock;
  assign axiDIO_reset = reset;
  assign axiDIO_io_axiIO_awready = io_dmaster_awready; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_wready = io_dmaster_wready; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_bvalid = io_dmaster_bvalid; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_arready = io_dmaster_arready; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_rvalid = io_dmaster_rvalid; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_rdata = io_dmaster_rdata; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_axiIO_rlast = io_dmaster_rlast; // @[ysyx_22041728.scala 256:21]
  assign axiDIO_io_cache_ar_valid_o = dCache_io_cacheOut_ar_valid_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_ar_addr_o = dCache_io_cacheOut_ar_addr_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_ar_len_o = dCache_io_cacheOut_ar_len_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_w_valid_o = dCache_io_cacheOut_w_valid_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_w_data_o = dCache_io_cacheOut_w_data_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_w_addr_o = dCache_io_cacheOut_w_addr_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_w_mask_o = dCache_io_cacheOut_w_mask_o; // @[ysyx_22041728.scala 48:18]
  assign axiDIO_io_cache_wsize = dCache_io_cacheOut_wsize; // @[ysyx_22041728.scala 48:18]
  assign imem_clock = clock;
  assign imem_io_memIO_cen = iCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 55:20]
  assign imem_io_memIO_wen = iCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 55:20]
  assign imem_io_memIO_wdata = iCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 55:20]
  assign imem_io_memIO_addr = iCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 55:20]
  assign imem_io_memIO_wmask = iCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 55:20]
  assign dmem_clock = clock;
  assign dmem_io_memIO_cen = dCache_io_SRAMIO_0_cen; // @[ysyx_22041728.scala 56:20]
  assign dmem_io_memIO_wen = dCache_io_SRAMIO_0_wen; // @[ysyx_22041728.scala 56:20]
  assign dmem_io_memIO_wdata = dCache_io_SRAMIO_0_wdata; // @[ysyx_22041728.scala 56:20]
  assign dmem_io_memIO_addr = dCache_io_SRAMIO_0_addr; // @[ysyx_22041728.scala 56:20]
  assign dmem_io_memIO_wmask = dCache_io_SRAMIO_0_wmask; // @[ysyx_22041728.scala 56:20]
  assign imem_1_clock = clock;
  assign imem_1_io_memIO_cen = iCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 55:20]
  assign imem_1_io_memIO_wen = iCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 55:20]
  assign imem_1_io_memIO_wdata = iCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 55:20]
  assign imem_1_io_memIO_addr = iCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 55:20]
  assign imem_1_io_memIO_wmask = iCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 55:20]
  assign dmem_1_clock = clock;
  assign dmem_1_io_memIO_cen = dCache_io_SRAMIO_1_cen; // @[ysyx_22041728.scala 56:20]
  assign dmem_1_io_memIO_wen = dCache_io_SRAMIO_1_wen; // @[ysyx_22041728.scala 56:20]
  assign dmem_1_io_memIO_wdata = dCache_io_SRAMIO_1_wdata; // @[ysyx_22041728.scala 56:20]
  assign dmem_1_io_memIO_addr = dCache_io_SRAMIO_1_addr; // @[ysyx_22041728.scala 56:20]
  assign dmem_1_io_memIO_wmask = dCache_io_SRAMIO_1_wmask; // @[ysyx_22041728.scala 56:20]
  assign imem_2_clock = clock;
  assign imem_2_io_memIO_cen = iCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 55:20]
  assign imem_2_io_memIO_wen = iCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 55:20]
  assign imem_2_io_memIO_wdata = iCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 55:20]
  assign imem_2_io_memIO_addr = iCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 55:20]
  assign imem_2_io_memIO_wmask = iCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 55:20]
  assign dmem_2_clock = clock;
  assign dmem_2_io_memIO_cen = dCache_io_SRAMIO_2_cen; // @[ysyx_22041728.scala 56:20]
  assign dmem_2_io_memIO_wen = dCache_io_SRAMIO_2_wen; // @[ysyx_22041728.scala 56:20]
  assign dmem_2_io_memIO_wdata = dCache_io_SRAMIO_2_wdata; // @[ysyx_22041728.scala 56:20]
  assign dmem_2_io_memIO_addr = dCache_io_SRAMIO_2_addr; // @[ysyx_22041728.scala 56:20]
  assign dmem_2_io_memIO_wmask = dCache_io_SRAMIO_2_wmask; // @[ysyx_22041728.scala 56:20]
  assign imem_3_clock = clock;
  assign imem_3_io_memIO_cen = iCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 55:20]
  assign imem_3_io_memIO_wen = iCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 55:20]
  assign imem_3_io_memIO_wdata = iCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 55:20]
  assign imem_3_io_memIO_addr = iCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 55:20]
  assign imem_3_io_memIO_wmask = iCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 55:20]
  assign dmem_3_clock = clock;
  assign dmem_3_io_memIO_cen = dCache_io_SRAMIO_3_cen; // @[ysyx_22041728.scala 56:20]
  assign dmem_3_io_memIO_wen = dCache_io_SRAMIO_3_wen; // @[ysyx_22041728.scala 56:20]
  assign dmem_3_io_memIO_wdata = dCache_io_SRAMIO_3_wdata; // @[ysyx_22041728.scala 56:20]
  assign dmem_3_io_memIO_addr = dCache_io_SRAMIO_3_addr; // @[ysyx_22041728.scala 56:20]
  assign dmem_3_io_memIO_wmask = dCache_io_SRAMIO_3_wmask; // @[ysyx_22041728.scala 56:20]
endmodule
